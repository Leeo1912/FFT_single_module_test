`timescale 1ns/1ps
module rom_4_rfft_data64
(
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic                     valid,
    input  logic [10:0]              addr_col1,
    input  logic [10:0]              addr_col2,
    output logic [63:0]              data_o_col1,
    output logic [63:0]              data_o_col2
);

    logic [63:0] coff[2047:0];

    assign coff[0   ] = 64'hffffa57effffa57e;
    assign coff[1   ] = 64'hffff89beffffcf04;
    assign coff[2   ] = 64'hffff9592ffffb8e3;
    assign coff[3   ] = 64'hffff8276ffffe707;
    assign coff[4   ] = 64'hffff8583ffffdad8;
    assign coff[5   ] = 64'hffff8f1dffffc3a9;
    assign coff[6   ] = 64'hffff9d0effffaecc;
    assign coff[7   ] = 64'hffff809efffff374;
    assign coff[8   ] = 64'hffff8163ffffed38;
    assign coff[9   ] = 64'hffff9930ffffb3c0;
    assign coff[10  ] = 64'hffff9236ffffbe32;
    assign coff[11  ] = 64'hffff83d6ffffe0e6;
    assign coff[12  ] = 64'hffff877bffffd4e1;
    assign coff[13  ] = 64'hffff8c4affffc946;
    assign coff[14  ] = 64'hffffa129ffffaa0a;
    assign coff[15  ] = 64'hffff8027fffff9b8;
    assign coff[16  ] = 64'hffff8059fffff695;
    assign coff[17  ] = 64'hffff9f14ffffac65;
    assign coff[18  ] = 64'hffff8dabffffc673;
    assign coff[19  ] = 64'hffff8676ffffd7d9;
    assign coff[20  ] = 64'hffff84a3ffffdddc;
    assign coff[21  ] = 64'hffff90a1ffffc0e9;
    assign coff[22  ] = 64'hffff9b17ffffb140;
    assign coff[23  ] = 64'hffff80f6fffff055;
    assign coff[24  ] = 64'hffff81e2ffffea1e;
    assign coff[25  ] = 64'hffff9759ffffb64c;
    assign coff[26  ] = 64'hffff93dcffffbb85;
    assign coff[27  ] = 64'hffff831cffffe3f4;
    assign coff[28  ] = 64'hffff8894ffffd1ef;
    assign coff[29  ] = 64'hffff8afbffffcc21;
    assign coff[30  ] = 64'hffffa34cffffa7bd;
    assign coff[31  ] = 64'hffff800afffffcdc;
    assign coff[32  ] = 64'hffff8016fffffb4a;
    assign coff[33  ] = 64'hffffa238ffffa8e2;
    assign coff[34  ] = 64'hffff8ba0ffffcab2;
    assign coff[35  ] = 64'hffff8805ffffd367;
    assign coff[36  ] = 64'hffff8377ffffe26d;
    assign coff[37  ] = 64'hffff9307ffffbcda;
    assign coff[38  ] = 64'hffff9843ffffb505;
    assign coff[39  ] = 64'hffff81a0ffffebab;
    assign coff[40  ] = 64'hffff812affffeec6;
    assign coff[41  ] = 64'hffff9a22ffffb27f;
    assign coff[42  ] = 64'hffff9169ffffbf8c;
    assign coff[43  ] = 64'hffff843affffdf61;
    assign coff[44  ] = 64'hffff86f6ffffd65c;
    assign coff[45  ] = 64'hffff8cf8ffffc7db;
    assign coff[46  ] = 64'hffffa01cffffab36;
    assign coff[47  ] = 64'hffff803efffff827;
    assign coff[48  ] = 64'hffff8079fffff505;
    assign coff[49  ] = 64'hffff9e0fffffad97;
    assign coff[50  ] = 64'hffff8e62ffffc50d;
    assign coff[51  ] = 64'hffff85faffffd958;
    assign coff[52  ] = 64'hffff8511ffffdc59;
    assign coff[53  ] = 64'hffff8fddffffc248;
    assign coff[54  ] = 64'hffff9c11ffffb005;
    assign coff[55  ] = 64'hffff80c8fffff1e4;
    assign coff[56  ] = 64'hffff822affffe892;
    assign coff[57  ] = 64'hffff9674ffffb796;
    assign coff[58  ] = 64'hffff94b5ffffba33;
    assign coff[59  ] = 64'hffff82c6ffffe57d;
    assign coff[60  ] = 64'hffff8927ffffd079;
    assign coff[61  ] = 64'hffff8a5affffcd92;
    assign coff[62  ] = 64'hffffa463ffffa69c;
    assign coff[63  ] = 64'hffff8002fffffe6e;
    assign coff[64  ] = 64'hffff8006fffffda5;
    assign coff[65  ] = 64'hffffa3d7ffffa72c;
    assign coff[66  ] = 64'hffff8aaaffffccd9;
    assign coff[67  ] = 64'hffff88ddffffd134;
    assign coff[68  ] = 64'hffff82f1ffffe4b9;
    assign coff[69  ] = 64'hffff9448ffffbadc;
    assign coff[70  ] = 64'hffff96e6ffffb6f1;
    assign coff[71  ] = 64'hffff8205ffffe958;
    assign coff[72  ] = 64'hffff80defffff11c;
    assign coff[73  ] = 64'hffff9b94ffffb0a2;
    assign coff[74  ] = 64'hffff903effffc198;
    assign coff[75  ] = 64'hffff84d9ffffdd1b;
    assign coff[76  ] = 64'hffff8637ffffd898;
    assign coff[77  ] = 64'hffff8e06ffffc5c0;
    assign coff[78  ] = 64'hffff9e91ffffacfd;
    assign coff[79  ] = 64'hffff8068fffff5cd;
    assign coff[80  ] = 64'hffff804bfffff75e;
    assign coff[81  ] = 64'hffff9f98ffffabcd;
    assign coff[82  ] = 64'hffff8d51ffffc727;
    assign coff[83  ] = 64'hffff86b6ffffd71b;
    assign coff[84  ] = 64'hffff846effffde9e;
    assign coff[85  ] = 64'hffff9105ffffc03a;
    assign coff[86  ] = 64'hffff9a9cffffb1df;
    assign coff[87  ] = 64'hffff8110ffffef8d;
    assign coff[88  ] = 64'hffff81c1ffffeae4;
    assign coff[89  ] = 64'hffff97ceffffb5a8;
    assign coff[90  ] = 64'hffff9371ffffbc2f;
    assign coff[91  ] = 64'hffff8349ffffe330;
    assign coff[92  ] = 64'hffff884cffffd2ab;
    assign coff[93  ] = 64'hffff8b4dffffcb69;
    assign coff[94  ] = 64'hffffa2c2ffffa84f;
    assign coff[95  ] = 64'hffff800ffffffc13;
    assign coff[96  ] = 64'hffff801efffffa81;
    assign coff[97  ] = 64'hffffa1b0ffffa976;
    assign coff[98  ] = 64'hffff8bf5ffffc9fc;
    assign coff[99  ] = 64'hffff87c0ffffd424;
    assign coff[100 ] = 64'hffff83a6ffffe1a9;
    assign coff[101 ] = 64'hffff929effffbd86;
    assign coff[102 ] = 64'hffff98b9ffffb462;
    assign coff[103 ] = 64'hffff8181ffffec71;
    assign coff[104 ] = 64'hffff8146ffffedff;
    assign coff[105 ] = 64'hffff99a9ffffb31f;
    assign coff[106 ] = 64'hffff91cfffffbedf;
    assign coff[107 ] = 64'hffff8407ffffe023;
    assign coff[108 ] = 64'hffff8738ffffd59e;
    assign coff[109 ] = 64'hffff8ca1ffffc890;
    assign coff[110 ] = 64'hffffa0a2ffffaaa0;
    assign coff[111 ] = 64'hffff8032fffff8ef;
    assign coff[112 ] = 64'hffff808bfffff43c;
    assign coff[113 ] = 64'hffff9d8effffae31;
    assign coff[114 ] = 64'hffff8ebfffffc45b;
    assign coff[115 ] = 64'hffff85beffffda18;
    assign coff[116 ] = 64'hffff8549ffffdb99;
    assign coff[117 ] = 64'hffff8f7dffffc2f8;
    assign coff[118 ] = 64'hffff9c8fffffaf68;
    assign coff[119 ] = 64'hffff80b2fffff2ac;
    assign coff[120 ] = 64'hffff824fffffe7cd;
    assign coff[121 ] = 64'hffff9603ffffb83c;
    assign coff[122 ] = 64'hffff9523ffffb98b;
    assign coff[123 ] = 64'hffff829dffffe642;
    assign coff[124 ] = 64'hffff8972ffffcfbe;
    assign coff[125 ] = 64'hffff8a0cffffce4b;
    assign coff[126 ] = 64'hffffa4f0ffffa60c;
    assign coff[127 ] = 64'hffff8001ffffff37;
    assign coff[128 ] = 64'hffff8001fffffed2;
    assign coff[129 ] = 64'hffffa4a9ffffa654;
    assign coff[130 ] = 64'hffff8a33ffffcdee;
    assign coff[131 ] = 64'hffff894cffffd01b;
    assign coff[132 ] = 64'hffff82b2ffffe5e0;
    assign coff[133 ] = 64'hffff94ecffffb9df;
    assign coff[134 ] = 64'hffff963bffffb7e9;
    assign coff[135 ] = 64'hffff823cffffe82f;
    assign coff[136 ] = 64'hffff80bdfffff248;
    assign coff[137 ] = 64'hffff9c50ffffafb6;
    assign coff[138 ] = 64'hffff8fadffffc2a0;
    assign coff[139 ] = 64'hffff852dffffdbf9;
    assign coff[140 ] = 64'hffff85dcffffd9b8;
    assign coff[141 ] = 64'hffff8e90ffffc4b4;
    assign coff[142 ] = 64'hffff9dceffffade4;
    assign coff[143 ] = 64'hffff8082fffff4a0;
    assign coff[144 ] = 64'hffff8038fffff88b;
    assign coff[145 ] = 64'hffffa05fffffaaeb;
    assign coff[146 ] = 64'hffff8cccffffc836;
    assign coff[147 ] = 64'hffff8717ffffd5fd;
    assign coff[148 ] = 64'hffff8421ffffdfc2;
    assign coff[149 ] = 64'hffff919cffffbf35;
    assign coff[150 ] = 64'hffff99e5ffffb2cf;
    assign coff[151 ] = 64'hffff8138ffffee62;
    assign coff[152 ] = 64'hffff8190ffffec0e;
    assign coff[153 ] = 64'hffff987effffb4b3;
    assign coff[154 ] = 64'hffff92d2ffffbd30;
    assign coff[155 ] = 64'hffff838effffe20b;
    assign coff[156 ] = 64'hffff87e2ffffd3c5;
    assign coff[157 ] = 64'hffff8bcaffffca57;
    assign coff[158 ] = 64'hffffa1f4ffffa92c;
    assign coff[159 ] = 64'hffff801afffffae5;
    assign coff[160 ] = 64'hffff8013fffffbae;
    assign coff[161 ] = 64'hffffa27dffffa899;
    assign coff[162 ] = 64'hffff8b77ffffcb0e;
    assign coff[163 ] = 64'hffff8828ffffd309;
    assign coff[164 ] = 64'hffff8360ffffe2cf;
    assign coff[165 ] = 64'hffff933cffffbc85;
    assign coff[166 ] = 64'hffff9808ffffb556;
    assign coff[167 ] = 64'hffff81b0ffffeb47;
    assign coff[168 ] = 64'hffff811dffffef2a;
    assign coff[169 ] = 64'hffff9a5fffffb22f;
    assign coff[170 ] = 64'hffff9137ffffbfe3;
    assign coff[171 ] = 64'hffff8454ffffdeff;
    assign coff[172 ] = 64'hffff86d6ffffd6bb;
    assign coff[173 ] = 64'hffff8d24ffffc781;
    assign coff[174 ] = 64'hffff9fdaffffab81;
    assign coff[175 ] = 64'hffff8044fffff7c2;
    assign coff[176 ] = 64'hffff8070fffff569;
    assign coff[177 ] = 64'hffff9e50ffffad4a;
    assign coff[178 ] = 64'hffff8e34ffffc566;
    assign coff[179 ] = 64'hffff8619ffffd8f8;
    assign coff[180 ] = 64'hffff84f5ffffdcba;
    assign coff[181 ] = 64'hffff900effffc1f0;
    assign coff[182 ] = 64'hffff9bd2ffffb053;
    assign coff[183 ] = 64'hffff80d3fffff180;
    assign coff[184 ] = 64'hffff8217ffffe8f5;
    assign coff[185 ] = 64'hffff96adffffb743;
    assign coff[186 ] = 64'hffff947effffba87;
    assign coff[187 ] = 64'hffff82dbffffe51b;
    assign coff[188 ] = 64'hffff8902ffffd0d6;
    assign coff[189 ] = 64'hffff8a82ffffcd35;
    assign coff[190 ] = 64'hffffa41dffffa6e4;
    assign coff[191 ] = 64'hffff8004fffffe09;
    assign coff[192 ] = 64'hffff8008fffffd40;
    assign coff[193 ] = 64'hffffa391ffffa774;
    assign coff[194 ] = 64'hffff8ad3ffffcc7d;
    assign coff[195 ] = 64'hffff88b8ffffd191;
    assign coff[196 ] = 64'hffff8306ffffe457;
    assign coff[197 ] = 64'hffff9412ffffbb30;
    assign coff[198 ] = 64'hffff9720ffffb69e;
    assign coff[199 ] = 64'hffff81f4ffffe9bb;
    assign coff[200 ] = 64'hffff80eafffff0b9;
    assign coff[201 ] = 64'hffff9b55ffffb0f1;
    assign coff[202 ] = 64'hffff9070ffffc140;
    assign coff[203 ] = 64'hffff84beffffdd7c;
    assign coff[204 ] = 64'hffff8656ffffd839;
    assign coff[205 ] = 64'hffff8dd8ffffc619;
    assign coff[206 ] = 64'hffff9ed2ffffacb1;
    assign coff[207 ] = 64'hffff8060fffff631;
    assign coff[208 ] = 64'hffff8052fffff6fa;
    assign coff[209 ] = 64'hffff9f56ffffac19;
    assign coff[210 ] = 64'hffff8d7effffc6cd;
    assign coff[211 ] = 64'hffff8696ffffd77a;
    assign coff[212 ] = 64'hffff8488ffffde3d;
    assign coff[213 ] = 64'hffff90d3ffffc091;
    assign coff[214 ] = 64'hffff9adaffffb18f;
    assign coff[215 ] = 64'hffff8103ffffeff1;
    assign coff[216 ] = 64'hffff81d1ffffea81;
    assign coff[217 ] = 64'hffff9793ffffb5fa;
    assign coff[218 ] = 64'hffff93a6ffffbbda;
    assign coff[219 ] = 64'hffff8332ffffe392;
    assign coff[220 ] = 64'hffff8870ffffd24d;
    assign coff[221 ] = 64'hffff8b24ffffcbc5;
    assign coff[222 ] = 64'hffffa307ffffa806;
    assign coff[223 ] = 64'hffff800cfffffc77;
    assign coff[224 ] = 64'hffff8023fffffa1d;
    assign coff[225 ] = 64'hffffa16cffffa9c0;
    assign coff[226 ] = 64'hffff8c1fffffc9a1;
    assign coff[227 ] = 64'hffff879dffffd482;
    assign coff[228 ] = 64'hffff83beffffe148;
    assign coff[229 ] = 64'hffff926affffbddc;
    assign coff[230 ] = 64'hffff98f5ffffb411;
    assign coff[231 ] = 64'hffff8172ffffecd5;
    assign coff[232 ] = 64'hffff8154ffffed9b;
    assign coff[233 ] = 64'hffff996dffffb36f;
    assign coff[234 ] = 64'hffff9202ffffbe88;
    assign coff[235 ] = 64'hffff83efffffe085;
    assign coff[236 ] = 64'hffff875affffd53f;
    assign coff[237 ] = 64'hffff8c75ffffc8eb;
    assign coff[238 ] = 64'hffffa0e5ffffaa55;
    assign coff[239 ] = 64'hffff802dfffff954;
    assign coff[240 ] = 64'hffff8094fffff3d8;
    assign coff[241 ] = 64'hffff9d4effffae7f;
    assign coff[242 ] = 64'hffff8eeeffffc402;
    assign coff[243 ] = 64'hffff85a0ffffda78;
    assign coff[244 ] = 64'hffff8566ffffdb38;
    assign coff[245 ] = 64'hffff8f4dffffc351;
    assign coff[246 ] = 64'hffff9cceffffaf1a;
    assign coff[247 ] = 64'hffff80a8fffff310;
    assign coff[248 ] = 64'hffff8262ffffe76a;
    assign coff[249 ] = 64'hffff95caffffb890;
    assign coff[250 ] = 64'hffff955bffffb937;
    assign coff[251 ] = 64'hffff8289ffffe6a5;
    assign coff[252 ] = 64'hffff8998ffffcf61;
    assign coff[253 ] = 64'hffff89e5ffffcea7;
    assign coff[254 ] = 64'hffffa537ffffa5c5;
    assign coff[255 ] = 64'hffff8000ffffff9b;
    assign coff[256 ] = 64'hffff8000ffffff69;
    assign coff[257 ] = 64'hffffa513ffffa5e8;
    assign coff[258 ] = 64'hffff89f8ffffce79;
    assign coff[259 ] = 64'hffff8985ffffcf90;
    assign coff[260 ] = 64'hffff8293ffffe673;
    assign coff[261 ] = 64'hffff953fffffb961;
    assign coff[262 ] = 64'hffff95e6ffffb866;
    assign coff[263 ] = 64'hffff8259ffffe79b;
    assign coff[264 ] = 64'hffff80adfffff2de;
    assign coff[265 ] = 64'hffff9cafffffaf41;
    assign coff[266 ] = 64'hffff8f65ffffc324;
    assign coff[267 ] = 64'hffff8558ffffdb68;
    assign coff[268 ] = 64'hffff85afffffda48;
    assign coff[269 ] = 64'hffff8ed6ffffc42e;
    assign coff[270 ] = 64'hffff9d6effffae58;
    assign coff[271 ] = 64'hffff808ffffff40a;
    assign coff[272 ] = 64'hffff802ffffff922;
    assign coff[273 ] = 64'hffffa0c4ffffaa7a;
    assign coff[274 ] = 64'hffff8c8bffffc8be;
    assign coff[275 ] = 64'hffff8749ffffd56f;
    assign coff[276 ] = 64'hffff83fbffffe054;
    assign coff[277 ] = 64'hffff91e9ffffbeb3;
    assign coff[278 ] = 64'hffff998bffffb347;
    assign coff[279 ] = 64'hffff814dffffedcd;
    assign coff[280 ] = 64'hffff8179ffffeca3;
    assign coff[281 ] = 64'hffff98d7ffffb439;
    assign coff[282 ] = 64'hffff9284ffffbdb1;
    assign coff[283 ] = 64'hffff83b2ffffe178;
    assign coff[284 ] = 64'hffff87afffffd453;
    assign coff[285 ] = 64'hffff8c0affffc9ce;
    assign coff[286 ] = 64'hffffa18effffa99b;
    assign coff[287 ] = 64'hffff8020fffffa4f;
    assign coff[288 ] = 64'hffff800efffffc45;
    assign coff[289 ] = 64'hffffa2e4ffffa82b;
    assign coff[290 ] = 64'hffff8b39ffffcb97;
    assign coff[291 ] = 64'hffff885effffd27c;
    assign coff[292 ] = 64'hffff833effffe361;
    assign coff[293 ] = 64'hffff938bffffbc05;
    assign coff[294 ] = 64'hffff97b0ffffb5d1;
    assign coff[295 ] = 64'hffff81c9ffffeab3;
    assign coff[296 ] = 64'hffff8109ffffefbf;
    assign coff[297 ] = 64'hffff9abbffffb1b7;
    assign coff[298 ] = 64'hffff90ecffffc066;
    assign coff[299 ] = 64'hffff847bffffde6e;
    assign coff[300 ] = 64'hffff86a5ffffd74a;
    assign coff[301 ] = 64'hffff8d67ffffc6fa;
    assign coff[302 ] = 64'hffff9f77ffffabf3;
    assign coff[303 ] = 64'hffff804efffff72c;
    assign coff[304 ] = 64'hffff8064fffff5ff;
    assign coff[305 ] = 64'hffff9eb2ffffacd7;
    assign coff[306 ] = 64'hffff8defffffc5ed;
    assign coff[307 ] = 64'hffff8647ffffd869;
    assign coff[308 ] = 64'hffff84ccffffdd4b;
    assign coff[309 ] = 64'hffff9057ffffc16c;
    assign coff[310 ] = 64'hffff9b75ffffb0c9;
    assign coff[311 ] = 64'hffff80e4fffff0eb;
    assign coff[312 ] = 64'hffff81fdffffe989;
    assign coff[313 ] = 64'hffff9703ffffb6c7;
    assign coff[314 ] = 64'hffff942dffffbb06;
    assign coff[315 ] = 64'hffff82fbffffe488;
    assign coff[316 ] = 64'hffff88caffffd162;
    assign coff[317 ] = 64'hffff8abeffffccab;
    assign coff[318 ] = 64'hffffa3b4ffffa750;
    assign coff[319 ] = 64'hffff8007fffffd73;
    assign coff[320 ] = 64'hffff8005fffffdd7;
    assign coff[321 ] = 64'hffffa3faffffa708;
    assign coff[322 ] = 64'hffff8a96ffffcd07;
    assign coff[323 ] = 64'hffff88efffffd105;
    assign coff[324 ] = 64'hffff82e6ffffe4ea;
    assign coff[325 ] = 64'hffff9463ffffbab1;
    assign coff[326 ] = 64'hffff96c9ffffb71a;
    assign coff[327 ] = 64'hffff820effffe926;
    assign coff[328 ] = 64'hffff80d9fffff14e;
    assign coff[329 ] = 64'hffff9bb3ffffb07b;
    assign coff[330 ] = 64'hffff9026ffffc1c4;
    assign coff[331 ] = 64'hffff84e7ffffdcea;
    assign coff[332 ] = 64'hffff8628ffffd8c8;
    assign coff[333 ] = 64'hffff8e1dffffc593;
    assign coff[334 ] = 64'hffff9e70ffffad24;
    assign coff[335 ] = 64'hffff806cfffff59b;
    assign coff[336 ] = 64'hffff8047fffff790;
    assign coff[337 ] = 64'hffff9fb9ffffaba7;
    assign coff[338 ] = 64'hffff8d3bffffc754;
    assign coff[339 ] = 64'hffff86c6ffffd6eb;
    assign coff[340 ] = 64'hffff8461ffffdecf;
    assign coff[341 ] = 64'hffff911effffc00f;
    assign coff[342 ] = 64'hffff9a7effffb207;
    assign coff[343 ] = 64'hffff8116ffffef5c;
    assign coff[344 ] = 64'hffff81b8ffffeb16;
    assign coff[345 ] = 64'hffff97ebffffb57f;
    assign coff[346 ] = 64'hffff9356ffffbc5a;
    assign coff[347 ] = 64'hffff8354ffffe2ff;
    assign coff[348 ] = 64'hffff883affffd2da;
    assign coff[349 ] = 64'hffff8b62ffffcb3c;
    assign coff[350 ] = 64'hffffa29fffffa874;
    assign coff[351 ] = 64'hffff8011fffffbe1;
    assign coff[352 ] = 64'hffff801cfffffab3;
    assign coff[353 ] = 64'hffffa1d2ffffa951;
    assign coff[354 ] = 64'hffff8bdfffffca29;
    assign coff[355 ] = 64'hffff87d1ffffd3f4;
    assign coff[356 ] = 64'hffff839affffe1da;
    assign coff[357 ] = 64'hffff92b8ffffbd5b;
    assign coff[358 ] = 64'hffff989cffffb48b;
    assign coff[359 ] = 64'hffff8188ffffec3f;
    assign coff[360 ] = 64'hffff813fffffee31;
    assign coff[361 ] = 64'hffff99c7ffffb2f7;
    assign coff[362 ] = 64'hffff91b6ffffbf0a;
    assign coff[363 ] = 64'hffff8414ffffdff2;
    assign coff[364 ] = 64'hffff8728ffffd5ce;
    assign coff[365 ] = 64'hffff8cb6ffffc863;
    assign coff[366 ] = 64'hffffa080ffffaac5;
    assign coff[367 ] = 64'hffff8035fffff8bd;
    assign coff[368 ] = 64'hffff8086fffff46e;
    assign coff[369 ] = 64'hffff9daeffffae0b;
    assign coff[370 ] = 64'hffff8ea8ffffc487;
    assign coff[371 ] = 64'hffff85cdffffd9e8;
    assign coff[372 ] = 64'hffff853bffffdbc9;
    assign coff[373 ] = 64'hffff8f95ffffc2cc;
    assign coff[374 ] = 64'hffff9c6fffffaf8f;
    assign coff[375 ] = 64'hffff80b7fffff27a;
    assign coff[376 ] = 64'hffff8246ffffe7fe;
    assign coff[377 ] = 64'hffff961fffffb813;
    assign coff[378 ] = 64'hffff9508ffffb9b5;
    assign coff[379 ] = 64'hffff82a8ffffe611;
    assign coff[380 ] = 64'hffff895fffffcfed;
    assign coff[381 ] = 64'hffff8a1fffffce1c;
    assign coff[382 ] = 64'hffffa4ccffffa630;
    assign coff[383 ] = 64'hffff8001ffffff05;
    assign coff[384 ] = 64'hffff8002fffffea0;
    assign coff[385 ] = 64'hffffa486ffffa678;
    assign coff[386 ] = 64'hffff8a47ffffcdc0;
    assign coff[387 ] = 64'hffff8939ffffd04a;
    assign coff[388 ] = 64'hffff82bcffffe5af;
    assign coff[389 ] = 64'hffff94d0ffffba09;
    assign coff[390 ] = 64'hffff9657ffffb7c0;
    assign coff[391 ] = 64'hffff8233ffffe861;
    assign coff[392 ] = 64'hffff80c2fffff216;
    assign coff[393 ] = 64'hffff9c30ffffafdd;
    assign coff[394 ] = 64'hffff8fc5ffffc274;
    assign coff[395 ] = 64'hffff851fffffdc29;
    assign coff[396 ] = 64'hffff85ebffffd988;
    assign coff[397 ] = 64'hffff8e79ffffc4e0;
    assign coff[398 ] = 64'hffff9defffffadbd;
    assign coff[399 ] = 64'hffff807dfffff4d3;
    assign coff[400 ] = 64'hffff803bfffff859;
    assign coff[401 ] = 64'hffffa03effffab10;
    assign coff[402 ] = 64'hffff8ce2ffffc809;
    assign coff[403 ] = 64'hffff8707ffffd62d;
    assign coff[404 ] = 64'hffff842dffffdf91;
    assign coff[405 ] = 64'hffff9183ffffbf61;
    assign coff[406 ] = 64'hffff9a04ffffb2a7;
    assign coff[407 ] = 64'hffff8131ffffee94;
    assign coff[408 ] = 64'hffff8198ffffebdc;
    assign coff[409 ] = 64'hffff9860ffffb4dc;
    assign coff[410 ] = 64'hffff92ecffffbd05;
    assign coff[411 ] = 64'hffff8382ffffe23c;
    assign coff[412 ] = 64'hffff87f4ffffd396;
    assign coff[413 ] = 64'hffff8bb5ffffca85;
    assign coff[414 ] = 64'hffffa216ffffa907;
    assign coff[415 ] = 64'hffff8018fffffb18;
    assign coff[416 ] = 64'hffff8014fffffb7c;
    assign coff[417 ] = 64'hffffa25bffffa8bd;
    assign coff[418 ] = 64'hffff8b8bffffcae0;
    assign coff[419 ] = 64'hffff8817ffffd338;
    assign coff[420 ] = 64'hffff836bffffe29e;
    assign coff[421 ] = 64'hffff9321ffffbcaf;
    assign coff[422 ] = 64'hffff9826ffffb52d;
    assign coff[423 ] = 64'hffff81a8ffffeb79;
    assign coff[424 ] = 64'hffff8123ffffeef8;
    assign coff[425 ] = 64'hffff9a40ffffb257;
    assign coff[426 ] = 64'hffff9150ffffbfb8;
    assign coff[427 ] = 64'hffff8447ffffdf30;
    assign coff[428 ] = 64'hffff86e6ffffd68c;
    assign coff[429 ] = 64'hffff8d0effffc7ae;
    assign coff[430 ] = 64'hffff9ffbffffab5c;
    assign coff[431 ] = 64'hffff8041fffff7f4;
    assign coff[432 ] = 64'hffff8075fffff537;
    assign coff[433 ] = 64'hffff9e2fffffad70;
    assign coff[434 ] = 64'hffff8e4bffffc53a;
    assign coff[435 ] = 64'hffff8609ffffd928;
    assign coff[436 ] = 64'hffff8503ffffdc8a;
    assign coff[437 ] = 64'hffff8ff5ffffc21c;
    assign coff[438 ] = 64'hffff9bf1ffffb02c;
    assign coff[439 ] = 64'hffff80cdfffff1b2;
    assign coff[440 ] = 64'hffff8220ffffe8c4;
    assign coff[441 ] = 64'hffff9690ffffb76d;
    assign coff[442 ] = 64'hffff949affffba5d;
    assign coff[443 ] = 64'hffff82d1ffffe54c;
    assign coff[444 ] = 64'hffff8914ffffd0a7;
    assign coff[445 ] = 64'hffff8a6effffcd63;
    assign coff[446 ] = 64'hffffa440ffffa6c0;
    assign coff[447 ] = 64'hffff8003fffffe3c;
    assign coff[448 ] = 64'hffff8009fffffd0e;
    assign coff[449 ] = 64'hffffa36fffffa799;
    assign coff[450 ] = 64'hffff8ae7ffffcc4f;
    assign coff[451 ] = 64'hffff88a6ffffd1c0;
    assign coff[452 ] = 64'hffff8311ffffe426;
    assign coff[453 ] = 64'hffff93f7ffffbb5b;
    assign coff[454 ] = 64'hffff973cffffb675;
    assign coff[455 ] = 64'hffff81ebffffe9ec;
    assign coff[456 ] = 64'hffff80f0fffff087;
    assign coff[457 ] = 64'hffff9b36ffffb118;
    assign coff[458 ] = 64'hffff9088ffffc114;
    assign coff[459 ] = 64'hffff84b0ffffddac;
    assign coff[460 ] = 64'hffff8666ffffd809;
    assign coff[461 ] = 64'hffff8dc1ffffc646;
    assign coff[462 ] = 64'hffff9ef3ffffac8b;
    assign coff[463 ] = 64'hffff805dfffff663;
    assign coff[464 ] = 64'hffff8055fffff6c8;
    assign coff[465 ] = 64'hffff9f35ffffac3f;
    assign coff[466 ] = 64'hffff8d94ffffc6a0;
    assign coff[467 ] = 64'hffff8686ffffd7aa;
    assign coff[468 ] = 64'hffff8496ffffde0d;
    assign coff[469 ] = 64'hffff90baffffc0bd;
    assign coff[470 ] = 64'hffff9af9ffffb168;
    assign coff[471 ] = 64'hffff80fdfffff023;
    assign coff[472 ] = 64'hffff81daffffea4f;
    assign coff[473 ] = 64'hffff9776ffffb623;
    assign coff[474 ] = 64'hffff93c1ffffbbb0;
    assign coff[475 ] = 64'hffff8327ffffe3c3;
    assign coff[476 ] = 64'hffff8882ffffd21e;
    assign coff[477 ] = 64'hffff8b10ffffcbf3;
    assign coff[478 ] = 64'hffffa329ffffa7e2;
    assign coff[479 ] = 64'hffff800bfffffcaa;
    assign coff[480 ] = 64'hffff8025fffff9ea;
    assign coff[481 ] = 64'hffffa14affffa9e5;
    assign coff[482 ] = 64'hffff8c35ffffc973;
    assign coff[483 ] = 64'hffff878cffffd4b1;
    assign coff[484 ] = 64'hffff83caffffe117;
    assign coff[485 ] = 64'hffff9250ffffbe07;
    assign coff[486 ] = 64'hffff9913ffffb3e9;
    assign coff[487 ] = 64'hffff816affffed06;
    assign coff[488 ] = 64'hffff815bffffed6a;
    assign coff[489 ] = 64'hffff994effffb398;
    assign coff[490 ] = 64'hffff921cffffbe5d;
    assign coff[491 ] = 64'hffff83e2ffffe0b5;
    assign coff[492 ] = 64'hffff876bffffd510;
    assign coff[493 ] = 64'hffff8c60ffffc918;
    assign coff[494 ] = 64'hffffa107ffffaa30;
    assign coff[495 ] = 64'hffff802afffff986;
    assign coff[496 ] = 64'hffff8099fffff3a6;
    assign coff[497 ] = 64'hffff9d2effffaea5;
    assign coff[498 ] = 64'hffff8f06ffffc3d6;
    assign coff[499 ] = 64'hffff8592ffffdaa8;
    assign coff[500 ] = 64'hffff8574ffffdb08;
    assign coff[501 ] = 64'hffff8f35ffffc37d;
    assign coff[502 ] = 64'hffff9ceeffffaef3;
    assign coff[503 ] = 64'hffff80a3fffff342;
    assign coff[504 ] = 64'hffff826cffffe739;
    assign coff[505 ] = 64'hffff95aeffffb8b9;
    assign coff[506 ] = 64'hffff9577ffffb90d;
    assign coff[507 ] = 64'hffff827fffffe6d6;
    assign coff[508 ] = 64'hffff89abffffcf33;
    assign coff[509 ] = 64'hffff89d2ffffced6;
    assign coff[510 ] = 64'hffffa55affffa5a1;
    assign coff[511 ] = 64'hffff8000ffffffce;
    assign coff[512 ] = 64'hffff8000ffffffb5;
    assign coff[513 ] = 64'hffffa548ffffa5b3;
    assign coff[514 ] = 64'hffff89dbffffcebf;
    assign coff[515 ] = 64'hffff89a2ffffcf4a;
    assign coff[516 ] = 64'hffff8284ffffe6bd;
    assign coff[517 ] = 64'hffff9569ffffb922;
    assign coff[518 ] = 64'hffff95bcffffb8a4;
    assign coff[519 ] = 64'hffff8267ffffe751;
    assign coff[520 ] = 64'hffff80a5fffff329;
    assign coff[521 ] = 64'hffff9cdeffffaf07;
    assign coff[522 ] = 64'hffff8f41ffffc367;
    assign coff[523 ] = 64'hffff856dffffdb20;
    assign coff[524 ] = 64'hffff8599ffffda90;
    assign coff[525 ] = 64'hffff8efaffffc3ec;
    assign coff[526 ] = 64'hffff9d3effffae92;
    assign coff[527 ] = 64'hffff8096fffff3bf;
    assign coff[528 ] = 64'hffff802bfffff96d;
    assign coff[529 ] = 64'hffffa0f6ffffaa42;
    assign coff[530 ] = 64'hffff8c6affffc902;
    assign coff[531 ] = 64'hffff8762ffffd528;
    assign coff[532 ] = 64'hffff83e8ffffe09d;
    assign coff[533 ] = 64'hffff920fffffbe73;
    assign coff[534 ] = 64'hffff995dffffb384;
    assign coff[535 ] = 64'hffff8158ffffed83;
    assign coff[536 ] = 64'hffff816effffeced;
    assign coff[537 ] = 64'hffff9904ffffb3fd;
    assign coff[538 ] = 64'hffff925dffffbdf1;
    assign coff[539 ] = 64'hffff83c4ffffe12f;
    assign coff[540 ] = 64'hffff8795ffffd49a;
    assign coff[541 ] = 64'hffff8c2affffc98a;
    assign coff[542 ] = 64'hffffa15bffffa9d3;
    assign coff[543 ] = 64'hffff8024fffffa03;
    assign coff[544 ] = 64'hffff800cfffffc90;
    assign coff[545 ] = 64'hffffa318ffffa7f4;
    assign coff[546 ] = 64'hffff8b1affffcbdc;
    assign coff[547 ] = 64'hffff8879ffffd235;
    assign coff[548 ] = 64'hffff832dffffe3ab;
    assign coff[549 ] = 64'hffff93b4ffffbbc5;
    assign coff[550 ] = 64'hffff9785ffffb60e;
    assign coff[551 ] = 64'hffff81d6ffffea68;
    assign coff[552 ] = 64'hffff8100fffff00a;
    assign coff[553 ] = 64'hffff9ae9ffffb17c;
    assign coff[554 ] = 64'hffff90c6ffffc0a7;
    assign coff[555 ] = 64'hffff848fffffde25;
    assign coff[556 ] = 64'hffff868effffd792;
    assign coff[557 ] = 64'hffff8d89ffffc6b7;
    assign coff[558 ] = 64'hffff9f45ffffac2c;
    assign coff[559 ] = 64'hffff8053fffff6e1;
    assign coff[560 ] = 64'hffff805efffff64a;
    assign coff[561 ] = 64'hffff9ee3ffffac9e;
    assign coff[562 ] = 64'hffff8dcdffffc630;
    assign coff[563 ] = 64'hffff865effffd821;
    assign coff[564 ] = 64'hffff84b7ffffdd94;
    assign coff[565 ] = 64'hffff907cffffc12a;
    assign coff[566 ] = 64'hffff9b46ffffb105;
    assign coff[567 ] = 64'hffff80edfffff0a0;
    assign coff[568 ] = 64'hffff81efffffe9d4;
    assign coff[569 ] = 64'hffff972effffb68a;
    assign coff[570 ] = 64'hffff9404ffffbb46;
    assign coff[571 ] = 64'hffff830cffffe43e;
    assign coff[572 ] = 64'hffff88afffffd1a9;
    assign coff[573 ] = 64'hffff8addffffcc66;
    assign coff[574 ] = 64'hffffa380ffffa787;
    assign coff[575 ] = 64'hffff8008fffffd27;
    assign coff[576 ] = 64'hffff8003fffffe22;
    assign coff[577 ] = 64'hffffa42effffa6d2;
    assign coff[578 ] = 64'hffff8a78ffffcd4c;
    assign coff[579 ] = 64'hffff890bffffd0bf;
    assign coff[580 ] = 64'hffff82d6ffffe534;
    assign coff[581 ] = 64'hffff948cffffba72;
    assign coff[582 ] = 64'hffff969fffffb758;
    assign coff[583 ] = 64'hffff821cffffe8dc;
    assign coff[584 ] = 64'hffff80d0fffff199;
    assign coff[585 ] = 64'hffff9be2ffffb040;
    assign coff[586 ] = 64'hffff9001ffffc206;
    assign coff[587 ] = 64'hffff84fcffffdca2;
    assign coff[588 ] = 64'hffff8611ffffd910;
    assign coff[589 ] = 64'hffff8e3fffffc550;
    assign coff[590 ] = 64'hffff9e40ffffad5d;
    assign coff[591 ] = 64'hffff8072fffff550;
    assign coff[592 ] = 64'hffff8042fffff7db;
    assign coff[593 ] = 64'hffff9feaffffab6f;
    assign coff[594 ] = 64'hffff8d19ffffc798;
    assign coff[595 ] = 64'hffff86deffffd6a4;
    assign coff[596 ] = 64'hffff844dffffdf18;
    assign coff[597 ] = 64'hffff9143ffffbfcd;
    assign coff[598 ] = 64'hffff9a50ffffb243;
    assign coff[599 ] = 64'hffff8120ffffef11;
    assign coff[600 ] = 64'hffff81acffffeb60;
    assign coff[601 ] = 64'hffff9817ffffb542;
    assign coff[602 ] = 64'hffff932effffbc9a;
    assign coff[603 ] = 64'hffff8365ffffe2b6;
    assign coff[604 ] = 64'hffff8820ffffd320;
    assign coff[605 ] = 64'hffff8b81ffffcaf7;
    assign coff[606 ] = 64'hffffa26cffffa8ab;
    assign coff[607 ] = 64'hffff8014fffffb95;
    assign coff[608 ] = 64'hffff8019fffffaff;
    assign coff[609 ] = 64'hffffa205ffffa919;
    assign coff[610 ] = 64'hffff8bc0ffffca6e;
    assign coff[611 ] = 64'hffff87ebffffd3ae;
    assign coff[612 ] = 64'hffff8388ffffe223;
    assign coff[613 ] = 64'hffff92dfffffbd1a;
    assign coff[614 ] = 64'hffff986fffffb4c8;
    assign coff[615 ] = 64'hffff8194ffffebf5;
    assign coff[616 ] = 64'hffff8134ffffee7b;
    assign coff[617 ] = 64'hffff99f4ffffb2bb;
    assign coff[618 ] = 64'hffff918fffffbf4b;
    assign coff[619 ] = 64'hffff8427ffffdfa9;
    assign coff[620 ] = 64'hffff870fffffd615;
    assign coff[621 ] = 64'hffff8cd7ffffc81f;
    assign coff[622 ] = 64'hffffa04effffaafe;
    assign coff[623 ] = 64'hffff8039fffff872;
    assign coff[624 ] = 64'hffff807ffffff4b9;
    assign coff[625 ] = 64'hffff9ddfffffadd1;
    assign coff[626 ] = 64'hffff8e85ffffc4ca;
    assign coff[627 ] = 64'hffff85e3ffffd9a0;
    assign coff[628 ] = 64'hffff8526ffffdc11;
    assign coff[629 ] = 64'hffff8fb9ffffc28a;
    assign coff[630 ] = 64'hffff9c40ffffafca;
    assign coff[631 ] = 64'hffff80bffffff22f;
    assign coff[632 ] = 64'hffff8237ffffe848;
    assign coff[633 ] = 64'hffff9649ffffb7d4;
    assign coff[634 ] = 64'hffff94deffffb9f4;
    assign coff[635 ] = 64'hffff82b7ffffe5c7;
    assign coff[636 ] = 64'hffff8943ffffd033;
    assign coff[637 ] = 64'hffff8a3dffffcdd7;
    assign coff[638 ] = 64'hffffa498ffffa666;
    assign coff[639 ] = 64'hffff8002fffffeb9;
    assign coff[640 ] = 64'hffff8001fffffeec;
    assign coff[641 ] = 64'hffffa4bbffffa642;
    assign coff[642 ] = 64'hffff8a29ffffce05;
    assign coff[643 ] = 64'hffff8956ffffd004;
    assign coff[644 ] = 64'hffff82adffffe5f8;
    assign coff[645 ] = 64'hffff94faffffb9ca;
    assign coff[646 ] = 64'hffff962dffffb7fe;
    assign coff[647 ] = 64'hffff8241ffffe817;
    assign coff[648 ] = 64'hffff80bafffff261;
    assign coff[649 ] = 64'hffff9c60ffffafa3;
    assign coff[650 ] = 64'hffff8fa1ffffc2b6;
    assign coff[651 ] = 64'hffff8534ffffdbe1;
    assign coff[652 ] = 64'hffff85d4ffffd9d0;
    assign coff[653 ] = 64'hffff8e9cffffc49e;
    assign coff[654 ] = 64'hffff9dbeffffadf7;
    assign coff[655 ] = 64'hffff8084fffff487;
    assign coff[656 ] = 64'hffff8036fffff8a4;
    assign coff[657 ] = 64'hffffa070ffffaad8;
    assign coff[658 ] = 64'hffff8cc1ffffc84c;
    assign coff[659 ] = 64'hffff871fffffd5e5;
    assign coff[660 ] = 64'hffff841affffdfda;
    assign coff[661 ] = 64'hffff91a9ffffbf20;
    assign coff[662 ] = 64'hffff99d6ffffb2e3;
    assign coff[663 ] = 64'hffff813bffffee4a;
    assign coff[664 ] = 64'hffff818cffffec27;
    assign coff[665 ] = 64'hffff988dffffb49f;
    assign coff[666 ] = 64'hffff92c5ffffbd45;
    assign coff[667 ] = 64'hffff8394ffffe1f2;
    assign coff[668 ] = 64'hffff87daffffd3dd;
    assign coff[669 ] = 64'hffff8bd5ffffca40;
    assign coff[670 ] = 64'hffffa1e3ffffa93e;
    assign coff[671 ] = 64'hffff801bfffffacc;
    assign coff[672 ] = 64'hffff8012fffffbc7;
    assign coff[673 ] = 64'hffffa28effffa886;
    assign coff[674 ] = 64'hffff8b6cffffcb25;
    assign coff[675 ] = 64'hffff8831ffffd2f1;
    assign coff[676 ] = 64'hffff835affffe2e7;
    assign coff[677 ] = 64'hffff9349ffffbc6f;
    assign coff[678 ] = 64'hffff97faffffb56b;
    assign coff[679 ] = 64'hffff81b4ffffeb2f;
    assign coff[680 ] = 64'hffff8119ffffef43;
    assign coff[681 ] = 64'hffff9a6effffb21b;
    assign coff[682 ] = 64'hffff912affffbff9;
    assign coff[683 ] = 64'hffff845affffdee7;
    assign coff[684 ] = 64'hffff86ceffffd6d3;
    assign coff[685 ] = 64'hffff8d30ffffc76b;
    assign coff[686 ] = 64'hffff9fc9ffffab94;
    assign coff[687 ] = 64'hffff8046fffff7a9;
    assign coff[688 ] = 64'hffff806efffff582;
    assign coff[689 ] = 64'hffff9e60ffffad37;
    assign coff[690 ] = 64'hffff8e28ffffc57d;
    assign coff[691 ] = 64'hffff8620ffffd8e0;
    assign coff[692 ] = 64'hffff84eeffffdcd2;
    assign coff[693 ] = 64'hffff901affffc1da;
    assign coff[694 ] = 64'hffff9bc2ffffb067;
    assign coff[695 ] = 64'hffff80d6fffff167;
    assign coff[696 ] = 64'hffff8213ffffe90e;
    assign coff[697 ] = 64'hffff96bbffffb72f;
    assign coff[698 ] = 64'hffff9471ffffba9c;
    assign coff[699 ] = 64'hffff82e1ffffe502;
    assign coff[700 ] = 64'hffff88f8ffffd0ed;
    assign coff[701 ] = 64'hffff8a8cffffcd1e;
    assign coff[702 ] = 64'hffffa40bffffa6f6;
    assign coff[703 ] = 64'hffff8004fffffdf0;
    assign coff[704 ] = 64'hffff8007fffffd59;
    assign coff[705 ] = 64'hffffa3a3ffffa762;
    assign coff[706 ] = 64'hffff8ac8ffffcc94;
    assign coff[707 ] = 64'hffff88c1ffffd17a;
    assign coff[708 ] = 64'hffff8301ffffe46f;
    assign coff[709 ] = 64'hffff941fffffbb1b;
    assign coff[710 ] = 64'hffff9711ffffb6b3;
    assign coff[711 ] = 64'hffff81f8ffffe9a2;
    assign coff[712 ] = 64'hffff80e7fffff0d2;
    assign coff[713 ] = 64'hffff9b65ffffb0dd;
    assign coff[714 ] = 64'hffff9063ffffc156;
    assign coff[715 ] = 64'hffff84c5ffffdd63;
    assign coff[716 ] = 64'hffff864fffffd851;
    assign coff[717 ] = 64'hffff8de4ffffc603;
    assign coff[718 ] = 64'hffff9ec2ffffacc4;
    assign coff[719 ] = 64'hffff8062fffff618;
    assign coff[720 ] = 64'hffff8050fffff713;
    assign coff[721 ] = 64'hffff9f66ffffac06;
    assign coff[722 ] = 64'hffff8d73ffffc6e3;
    assign coff[723 ] = 64'hffff869effffd762;
    assign coff[724 ] = 64'hffff8482ffffde56;
    assign coff[725 ] = 64'hffff90dfffffc07b;
    assign coff[726 ] = 64'hffff9acaffffb1a3;
    assign coff[727 ] = 64'hffff8106ffffefd8;
    assign coff[728 ] = 64'hffff81cdffffea9a;
    assign coff[729 ] = 64'hffff97a2ffffb5e5;
    assign coff[730 ] = 64'hffff9399ffffbbef;
    assign coff[731 ] = 64'hffff8338ffffe37a;
    assign coff[732 ] = 64'hffff8867ffffd264;
    assign coff[733 ] = 64'hffff8b2effffcbae;
    assign coff[734 ] = 64'hffffa2f5ffffa818;
    assign coff[735 ] = 64'hffff800dfffffc5e;
    assign coff[736 ] = 64'hffff8022fffffa36;
    assign coff[737 ] = 64'hffffa17dffffa9ad;
    assign coff[738 ] = 64'hffff8c15ffffc9b8;
    assign coff[739 ] = 64'hffff87a6ffffd46b;
    assign coff[740 ] = 64'hffff83b8ffffe160;
    assign coff[741 ] = 64'hffff9277ffffbdc6;
    assign coff[742 ] = 64'hffff98e6ffffb425;
    assign coff[743 ] = 64'hffff8175ffffecbc;
    assign coff[744 ] = 64'hffff8150ffffedb4;
    assign coff[745 ] = 64'hffff997cffffb35b;
    assign coff[746 ] = 64'hffff91f6ffffbe9e;
    assign coff[747 ] = 64'hffff83f5ffffe06c;
    assign coff[748 ] = 64'hffff8751ffffd557;
    assign coff[749 ] = 64'hffff8c80ffffc8d4;
    assign coff[750 ] = 64'hffffa0d4ffffaa68;
    assign coff[751 ] = 64'hffff802efffff93b;
    assign coff[752 ] = 64'hffff8092fffff3f1;
    assign coff[753 ] = 64'hffff9d5effffae6b;
    assign coff[754 ] = 64'hffff8ee2ffffc418;
    assign coff[755 ] = 64'hffff85a8ffffda60;
    assign coff[756 ] = 64'hffff855fffffdb50;
    assign coff[757 ] = 64'hffff8f59ffffc33b;
    assign coff[758 ] = 64'hffff9cbeffffaf2d;
    assign coff[759 ] = 64'hffff80aafffff2f7;
    assign coff[760 ] = 64'hffff825dffffe783;
    assign coff[761 ] = 64'hffff95d8ffffb87b;
    assign coff[762 ] = 64'hffff954dffffb94c;
    assign coff[763 ] = 64'hffff828effffe68c;
    assign coff[764 ] = 64'hffff898effffcf78;
    assign coff[765 ] = 64'hffff89efffffce90;
    assign coff[766 ] = 64'hffffa525ffffa5d7;
    assign coff[767 ] = 64'hffff8000ffffff82;
    assign coff[768 ] = 64'hffff8000ffffff50;
    assign coff[769 ] = 64'hffffa501ffffa5fa;
    assign coff[770 ] = 64'hffff8a02ffffce62;
    assign coff[771 ] = 64'hffff897bffffcfa7;
    assign coff[772 ] = 64'hffff8298ffffe65b;
    assign coff[773 ] = 64'hffff9531ffffb976;
    assign coff[774 ] = 64'hffff95f5ffffb851;
    assign coff[775 ] = 64'hffff8254ffffe7b4;
    assign coff[776 ] = 64'hffff80b0fffff2c5;
    assign coff[777 ] = 64'hffff9c9fffffaf54;
    assign coff[778 ] = 64'hffff8f71ffffc30e;
    assign coff[779 ] = 64'hffff8550ffffdb80;
    assign coff[780 ] = 64'hffff85b7ffffda30;
    assign coff[781 ] = 64'hffff8ecbffffc445;
    assign coff[782 ] = 64'hffff9d7effffae45;
    assign coff[783 ] = 64'hffff808dfffff423;
    assign coff[784 ] = 64'hffff8031fffff908;
    assign coff[785 ] = 64'hffffa0b3ffffaa8d;
    assign coff[786 ] = 64'hffff8c96ffffc8a7;
    assign coff[787 ] = 64'hffff8741ffffd587;
    assign coff[788 ] = 64'hffff8401ffffe03b;
    assign coff[789 ] = 64'hffff91dcffffbec9;
    assign coff[790 ] = 64'hffff999affffb333;
    assign coff[791 ] = 64'hffff8149ffffede6;
    assign coff[792 ] = 64'hffff817dffffec8a;
    assign coff[793 ] = 64'hffff98c8ffffb44e;
    assign coff[794 ] = 64'hffff9291ffffbd9b;
    assign coff[795 ] = 64'hffff83acffffe191;
    assign coff[796 ] = 64'hffff87b7ffffd43b;
    assign coff[797 ] = 64'hffff8bffffffc9e5;
    assign coff[798 ] = 64'hffffa19fffffa988;
    assign coff[799 ] = 64'hffff801ffffffa68;
    assign coff[800 ] = 64'hffff800ffffffc2c;
    assign coff[801 ] = 64'hffffa2d3ffffa83d;
    assign coff[802 ] = 64'hffff8b43ffffcb80;
    assign coff[803 ] = 64'hffff8855ffffd293;
    assign coff[804 ] = 64'hffff8343ffffe349;
    assign coff[805 ] = 64'hffff937effffbc1a;
    assign coff[806 ] = 64'hffff97bfffffb5bc;
    assign coff[807 ] = 64'hffff81c5ffffeacb;
    assign coff[808 ] = 64'hffff810cffffefa6;
    assign coff[809 ] = 64'hffff9aacffffb1cb;
    assign coff[810 ] = 64'hffff90f8ffffc050;
    assign coff[811 ] = 64'hffff8475ffffde86;
    assign coff[812 ] = 64'hffff86adffffd732;
    assign coff[813 ] = 64'hffff8d5cffffc710;
    assign coff[814 ] = 64'hffff9f87ffffabe0;
    assign coff[815 ] = 64'hffff804cfffff745;
    assign coff[816 ] = 64'hffff8066fffff5e6;
    assign coff[817 ] = 64'hffff9ea1ffffacea;
    assign coff[818 ] = 64'hffff8dfaffffc5d6;
    assign coff[819 ] = 64'hffff863fffffd880;
    assign coff[820 ] = 64'hffff84d2ffffdd33;
    assign coff[821 ] = 64'hffff904bffffc182;
    assign coff[822 ] = 64'hffff9b84ffffb0b6;
    assign coff[823 ] = 64'hffff80e1fffff104;
    assign coff[824 ] = 64'hffff8201ffffe971;
    assign coff[825 ] = 64'hffff96f4ffffb6dc;
    assign coff[826 ] = 64'hffff943affffbaf1;
    assign coff[827 ] = 64'hffff82f6ffffe4a0;
    assign coff[828 ] = 64'hffff88d3ffffd14b;
    assign coff[829 ] = 64'hffff8ab4ffffccc2;
    assign coff[830 ] = 64'hffffa3c6ffffa73e;
    assign coff[831 ] = 64'hffff8006fffffd8c;
    assign coff[832 ] = 64'hffff8005fffffdbe;
    assign coff[833 ] = 64'hffffa3e8ffffa71a;
    assign coff[834 ] = 64'hffff8aa0ffffccf0;
    assign coff[835 ] = 64'hffff88e6ffffd11c;
    assign coff[836 ] = 64'hffff82ebffffe4d1;
    assign coff[837 ] = 64'hffff9456ffffbac7;
    assign coff[838 ] = 64'hffff96d8ffffb705;
    assign coff[839 ] = 64'hffff820affffe93f;
    assign coff[840 ] = 64'hffff80dcfffff135;
    assign coff[841 ] = 64'hffff9ba3ffffb08e;
    assign coff[842 ] = 64'hffff9032ffffc1ae;
    assign coff[843 ] = 64'hffff84e0ffffdd03;
    assign coff[844 ] = 64'hffff8630ffffd8b0;
    assign coff[845 ] = 64'hffff8e11ffffc5a9;
    assign coff[846 ] = 64'hffff9e81ffffad11;
    assign coff[847 ] = 64'hffff806afffff5b4;
    assign coff[848 ] = 64'hffff8049fffff777;
    assign coff[849 ] = 64'hffff9fa8ffffabba;
    assign coff[850 ] = 64'hffff8d46ffffc73e;
    assign coff[851 ] = 64'hffff86beffffd703;
    assign coff[852 ] = 64'hffff8467ffffdeb7;
    assign coff[853 ] = 64'hffff9111ffffc024;
    assign coff[854 ] = 64'hffff9a8dffffb1f3;
    assign coff[855 ] = 64'hffff8113ffffef74;
    assign coff[856 ] = 64'hffff81bdffffeafd;
    assign coff[857 ] = 64'hffff97dcffffb593;
    assign coff[858 ] = 64'hffff9363ffffbc45;
    assign coff[859 ] = 64'hffff834fffffe318;
    assign coff[860 ] = 64'hffff8843ffffd2c2;
    assign coff[861 ] = 64'hffff8b58ffffcb53;
    assign coff[862 ] = 64'hffffa2b0ffffa861;
    assign coff[863 ] = 64'hffff8010fffffbfa;
    assign coff[864 ] = 64'hffff801dfffffa9a;
    assign coff[865 ] = 64'hffffa1c1ffffa963;
    assign coff[866 ] = 64'hffff8beaffffca13;
    assign coff[867 ] = 64'hffff87c8ffffd40c;
    assign coff[868 ] = 64'hffff83a0ffffe1c2;
    assign coff[869 ] = 64'hffff92abffffbd70;
    assign coff[870 ] = 64'hffff98aaffffb476;
    assign coff[871 ] = 64'hffff8185ffffec58;
    assign coff[872 ] = 64'hffff8142ffffee18;
    assign coff[873 ] = 64'hffff99b8ffffb30b;
    assign coff[874 ] = 64'hffff91c2ffffbef4;
    assign coff[875 ] = 64'hffff840effffe00b;
    assign coff[876 ] = 64'hffff8730ffffd5b6;
    assign coff[877 ] = 64'hffff8cabffffc87a;
    assign coff[878 ] = 64'hffffa091ffffaab2;
    assign coff[879 ] = 64'hffff8033fffff8d6;
    assign coff[880 ] = 64'hffff8088fffff455;
    assign coff[881 ] = 64'hffff9d9effffae1e;
    assign coff[882 ] = 64'hffff8eb3ffffc471;
    assign coff[883 ] = 64'hffff85c5ffffda00;
    assign coff[884 ] = 64'hffff8542ffffdbb1;
    assign coff[885 ] = 64'hffff8f89ffffc2e2;
    assign coff[886 ] = 64'hffff9c7fffffaf7c;
    assign coff[887 ] = 64'hffff80b5fffff293;
    assign coff[888 ] = 64'hffff824affffe7e5;
    assign coff[889 ] = 64'hffff9611ffffb827;
    assign coff[890 ] = 64'hffff9515ffffb9a0;
    assign coff[891 ] = 64'hffff82a3ffffe62a;
    assign coff[892 ] = 64'hffff8968ffffcfd6;
    assign coff[893 ] = 64'hffff8a16ffffce34;
    assign coff[894 ] = 64'hffffa4deffffa61e;
    assign coff[895 ] = 64'hffff8001ffffff1e;
    assign coff[896 ] = 64'hffff8002fffffe87;
    assign coff[897 ] = 64'hffffa474ffffa68a;
    assign coff[898 ] = 64'hffff8a51ffffcda9;
    assign coff[899 ] = 64'hffff8930ffffd061;
    assign coff[900 ] = 64'hffff82c1ffffe596;
    assign coff[901 ] = 64'hffff94c3ffffba1e;
    assign coff[902 ] = 64'hffff9666ffffb7ab;
    assign coff[903 ] = 64'hffff822effffe879;
    assign coff[904 ] = 64'hffff80c5fffff1fd;
    assign coff[905 ] = 64'hffff9c21ffffaff1;
    assign coff[906 ] = 64'hffff8fd1ffffc25e;
    assign coff[907 ] = 64'hffff8518ffffdc41;
    assign coff[908 ] = 64'hffff85f2ffffd970;
    assign coff[909 ] = 64'hffff8e6dffffc4f7;
    assign coff[910 ] = 64'hffff9dffffffadaa;
    assign coff[911 ] = 64'hffff807bfffff4ec;
    assign coff[912 ] = 64'hffff803cfffff840;
    assign coff[913 ] = 64'hffffa02dffffab23;
    assign coff[914 ] = 64'hffff8cedffffc7f2;
    assign coff[915 ] = 64'hffff86ffffffd644;
    assign coff[916 ] = 64'hffff8434ffffdf79;
    assign coff[917 ] = 64'hffff9176ffffbf76;
    assign coff[918 ] = 64'hffff9a13ffffb293;
    assign coff[919 ] = 64'hffff812dffffeead;
    assign coff[920 ] = 64'hffff819cffffebc3;
    assign coff[921 ] = 64'hffff9852ffffb4f0;
    assign coff[922 ] = 64'hffff92faffffbcf0;
    assign coff[923 ] = 64'hffff837dffffe254;
    assign coff[924 ] = 64'hffff87fdffffd37f;
    assign coff[925 ] = 64'hffff8babffffca9c;
    assign coff[926 ] = 64'hffffa227ffffa8f4;
    assign coff[927 ] = 64'hffff8017fffffb31;
    assign coff[928 ] = 64'hffff8015fffffb63;
    assign coff[929 ] = 64'hffffa249ffffa8d0;
    assign coff[930 ] = 64'hffff8b96ffffcac9;
    assign coff[931 ] = 64'hffff880effffd34f;
    assign coff[932 ] = 64'hffff8371ffffe285;
    assign coff[933 ] = 64'hffff9314ffffbcc5;
    assign coff[934 ] = 64'hffff9834ffffb519;
    assign coff[935 ] = 64'hffff81a4ffffeb92;
    assign coff[936 ] = 64'hffff8127ffffeedf;
    assign coff[937 ] = 64'hffff9a31ffffb26b;
    assign coff[938 ] = 64'hffff915dffffbfa2;
    assign coff[939 ] = 64'hffff8441ffffdf48;
    assign coff[940 ] = 64'hffff86eeffffd674;
    assign coff[941 ] = 64'hffff8d03ffffc7c5;
    assign coff[942 ] = 64'hffffa00cffffab49;
    assign coff[943 ] = 64'hffff803ffffff80e;
    assign coff[944 ] = 64'hffff8077fffff51e;
    assign coff[945 ] = 64'hffff9e1fffffad84;
    assign coff[946 ] = 64'hffff8e56ffffc523;
    assign coff[947 ] = 64'hffff8602ffffd940;
    assign coff[948 ] = 64'hffff850affffdc72;
    assign coff[949 ] = 64'hffff8fe9ffffc232;
    assign coff[950 ] = 64'hffff9c01ffffb018;
    assign coff[951 ] = 64'hffff80cafffff1cb;
    assign coff[952 ] = 64'hffff8225ffffe8ab;
    assign coff[953 ] = 64'hffff9682ffffb781;
    assign coff[954 ] = 64'hffff94a7ffffba48;
    assign coff[955 ] = 64'hffff82ccffffe565;
    assign coff[956 ] = 64'hffff891dffffd090;
    assign coff[957 ] = 64'hffff8a64ffffcd7b;
    assign coff[958 ] = 64'hffffa451ffffa6ae;
    assign coff[959 ] = 64'hffff8003fffffe55;
    assign coff[960 ] = 64'hffff8009fffffcf5;
    assign coff[961 ] = 64'hffffa35dffffa7ab;
    assign coff[962 ] = 64'hffff8af1ffffcc38;
    assign coff[963 ] = 64'hffff889dffffd1d8;
    assign coff[964 ] = 64'hffff8317ffffe40d;
    assign coff[965 ] = 64'hffff93e9ffffbb70;
    assign coff[966 ] = 64'hffff974bffffb660;
    assign coff[967 ] = 64'hffff81e7ffffea05;
    assign coff[968 ] = 64'hffff80f3fffff06e;
    assign coff[969 ] = 64'hffff9b27ffffb12c;
    assign coff[970 ] = 64'hffff9095ffffc0ff;
    assign coff[971 ] = 64'hffff84aaffffddc4;
    assign coff[972 ] = 64'hffff866effffd7f1;
    assign coff[973 ] = 64'hffff8db6ffffc65d;
    assign coff[974 ] = 64'hffff9f03ffffac78;
    assign coff[975 ] = 64'hffff805bfffff67c;
    assign coff[976 ] = 64'hffff8057fffff6af;
    assign coff[977 ] = 64'hffff9f24ffffac52;
    assign coff[978 ] = 64'hffff8da0ffffc68a;
    assign coff[979 ] = 64'hffff867effffd7c1;
    assign coff[980 ] = 64'hffff849cffffddf5;
    assign coff[981 ] = 64'hffff90adffffc0d3;
    assign coff[982 ] = 64'hffff9b08ffffb154;
    assign coff[983 ] = 64'hffff80fafffff03c;
    assign coff[984 ] = 64'hffff81deffffea37;
    assign coff[985 ] = 64'hffff9768ffffb637;
    assign coff[986 ] = 64'hffff93ceffffbb9a;
    assign coff[987 ] = 64'hffff8322ffffe3dc;
    assign coff[988 ] = 64'hffff888bffffd206;
    assign coff[989 ] = 64'hffff8b05ffffcc0a;
    assign coff[990 ] = 64'hffffa33bffffa7cf;
    assign coff[991 ] = 64'hffff800afffffcc3;
    assign coff[992 ] = 64'hffff8026fffff9d1;
    assign coff[993 ] = 64'hffffa139ffffa9f8;
    assign coff[994 ] = 64'hffff8c3fffffc95d;
    assign coff[995 ] = 64'hffff8784ffffd4c9;
    assign coff[996 ] = 64'hffff83d0ffffe0fe;
    assign coff[997 ] = 64'hffff9243ffffbe1c;
    assign coff[998 ] = 64'hffff9922ffffb3d4;
    assign coff[999 ] = 64'hffff8166ffffed1f;
    assign coff[1000] = 64'hffff815fffffed51;
    assign coff[1001] = 64'hffff993fffffb3ac;
    assign coff[1002] = 64'hffff9229ffffbe47;
    assign coff[1003] = 64'hffff83dcffffe0ce;
    assign coff[1004] = 64'hffff8773ffffd4f8;
    assign coff[1005] = 64'hffff8c55ffffc92f;
    assign coff[1006] = 64'hffffa118ffffaa1d;
    assign coff[1007] = 64'hffff8029fffff99f;
    assign coff[1008] = 64'hffff809bfffff38d;
    assign coff[1009] = 64'hffff9d1effffaeb9;
    assign coff[1010] = 64'hffff8f11ffffc3bf;
    assign coff[1011] = 64'hffff858affffdac0;
    assign coff[1012] = 64'hffff857cffffdaf0;
    assign coff[1013] = 64'hffff8f29ffffc393;
    assign coff[1014] = 64'hffff9cfeffffaee0;
    assign coff[1015] = 64'hffff80a0fffff35b;
    assign coff[1016] = 64'hffff8271ffffe720;
    assign coff[1017] = 64'hffff95a0ffffb8ce;
    assign coff[1018] = 64'hffff9584ffffb8f8;
    assign coff[1019] = 64'hffff827bffffe6ef;
    assign coff[1020] = 64'hffff89b5ffffcf1b;
    assign coff[1021] = 64'hffff89c8ffffceed;
    assign coff[1022] = 64'hffffa56cffffa58f;
    assign coff[1023] = 64'hffff8000ffffffe7;
    assign coff[1024] = 64'hffff8000ffffffda;
    assign coff[1025] = 64'hffffa563ffffa598;
    assign coff[1026] = 64'hffff89cdffffcee1;
    assign coff[1027] = 64'hffff89b0ffffcf27;
    assign coff[1028] = 64'hffff827dffffe6e2;
    assign coff[1029] = 64'hffff957dffffb902;
    assign coff[1030] = 64'hffff95a7ffffb8c4;
    assign coff[1031] = 64'hffff826effffe72c;
    assign coff[1032] = 64'hffff80a2fffff34f;
    assign coff[1033] = 64'hffff9cf6ffffaee9;
    assign coff[1034] = 64'hffff8f2fffffc388;
    assign coff[1035] = 64'hffff8578ffffdafc;
    assign coff[1036] = 64'hffff858effffdab4;
    assign coff[1037] = 64'hffff8f0bffffc3cb;
    assign coff[1038] = 64'hffff9d26ffffaeaf;
    assign coff[1039] = 64'hffff809afffff39a;
    assign coff[1040] = 64'hffff8029fffff992;
    assign coff[1041] = 64'hffffa10fffffaa26;
    assign coff[1042] = 64'hffff8c5affffc924;
    assign coff[1043] = 64'hffff876fffffd504;
    assign coff[1044] = 64'hffff83dfffffe0c1;
    assign coff[1045] = 64'hffff9223ffffbe52;
    assign coff[1046] = 64'hffff9947ffffb3a2;
    assign coff[1047] = 64'hffff815dffffed5d;
    assign coff[1048] = 64'hffff8168ffffed13;
    assign coff[1049] = 64'hffff991affffb3de;
    assign coff[1050] = 64'hffff9249ffffbe12;
    assign coff[1051] = 64'hffff83cdffffe10b;
    assign coff[1052] = 64'hffff8788ffffd4bd;
    assign coff[1053] = 64'hffff8c3affffc968;
    assign coff[1054] = 64'hffffa142ffffa9ee;
    assign coff[1055] = 64'hffff8026fffff9de;
    assign coff[1056] = 64'hffff800bfffffcb6;
    assign coff[1057] = 64'hffffa332ffffa7d8;
    assign coff[1058] = 64'hffff8b0affffcbff;
    assign coff[1059] = 64'hffff8886ffffd212;
    assign coff[1060] = 64'hffff8324ffffe3d0;
    assign coff[1061] = 64'hffff93c8ffffbba5;
    assign coff[1062] = 64'hffff976fffffb62d;
    assign coff[1063] = 64'hffff81dcffffea43;
    assign coff[1064] = 64'hffff80fbfffff02f;
    assign coff[1065] = 64'hffff9b00ffffb15e;
    assign coff[1066] = 64'hffff90b4ffffc0c8;
    assign coff[1067] = 64'hffff8499ffffde01;
    assign coff[1068] = 64'hffff8682ffffd7b5;
    assign coff[1069] = 64'hffff8d9affffc695;
    assign coff[1070] = 64'hffff9f2cffffac48;
    assign coff[1071] = 64'hffff8056fffff6bb;
    assign coff[1072] = 64'hffff805cfffff670;
    assign coff[1073] = 64'hffff9efbffffac81;
    assign coff[1074] = 64'hffff8dbcffffc651;
    assign coff[1075] = 64'hffff866affffd7fd;
    assign coff[1076] = 64'hffff84adffffddb8;
    assign coff[1077] = 64'hffff908effffc10a;
    assign coff[1078] = 64'hffff9b2fffffb122;
    assign coff[1079] = 64'hffff80f2fffff07a;
    assign coff[1080] = 64'hffff81e9ffffe9f9;
    assign coff[1081] = 64'hffff9744ffffb66b;
    assign coff[1082] = 64'hffff93f0ffffbb65;
    assign coff[1083] = 64'hffff8314ffffe419;
    assign coff[1084] = 64'hffff88a1ffffd1cc;
    assign coff[1085] = 64'hffff8aecffffcc44;
    assign coff[1086] = 64'hffffa366ffffa7a2;
    assign coff[1087] = 64'hffff8009fffffd02;
    assign coff[1088] = 64'hffff8003fffffe48;
    assign coff[1089] = 64'hffffa449ffffa6b7;
    assign coff[1090] = 64'hffff8a69ffffcd6f;
    assign coff[1091] = 64'hffff8919ffffd09c;
    assign coff[1092] = 64'hffff82ceffffe558;
    assign coff[1093] = 64'hffff94a1ffffba52;
    assign coff[1094] = 64'hffff9689ffffb777;
    assign coff[1095] = 64'hffff8223ffffe8b7;
    assign coff[1096] = 64'hffff80ccfffff1bf;
    assign coff[1097] = 64'hffff9bf9ffffb022;
    assign coff[1098] = 64'hffff8fefffffc227;
    assign coff[1099] = 64'hffff8506ffffdc7e;
    assign coff[1100] = 64'hffff8605ffffd934;
    assign coff[1101] = 64'hffff8e50ffffc52f;
    assign coff[1102] = 64'hffff9e27ffffad7a;
    assign coff[1103] = 64'hffff8076fffff52a;
    assign coff[1104] = 64'hffff8040fffff801;
    assign coff[1105] = 64'hffffa003ffffab52;
    assign coff[1106] = 64'hffff8d09ffffc7ba;
    assign coff[1107] = 64'hffff86eaffffd680;
    assign coff[1108] = 64'hffff8444ffffdf3c;
    assign coff[1109] = 64'hffff9156ffffbfad;
    assign coff[1110] = 64'hffff9a39ffffb261;
    assign coff[1111] = 64'hffff8125ffffeeeb;
    assign coff[1112] = 64'hffff81a6ffffeb85;
    assign coff[1113] = 64'hffff982dffffb523;
    assign coff[1114] = 64'hffff931bffffbcba;
    assign coff[1115] = 64'hffff836effffe291;
    assign coff[1116] = 64'hffff8812ffffd344;
    assign coff[1117] = 64'hffff8b91ffffcad5;
    assign coff[1118] = 64'hffffa252ffffa8c6;
    assign coff[1119] = 64'hffff8015fffffb70;
    assign coff[1120] = 64'hffff8018fffffb24;
    assign coff[1121] = 64'hffffa21fffffa8fe;
    assign coff[1122] = 64'hffff8bb0ffffca90;
    assign coff[1123] = 64'hffff87f8ffffd38a;
    assign coff[1124] = 64'hffff837fffffe248;
    assign coff[1125] = 64'hffff92f3ffffbcfa;
    assign coff[1126] = 64'hffff9859ffffb4e6;
    assign coff[1127] = 64'hffff819affffebd0;
    assign coff[1128] = 64'hffff812fffffeea1;
    assign coff[1129] = 64'hffff9a0bffffb29d;
    assign coff[1130] = 64'hffff917cffffbf6b;
    assign coff[1131] = 64'hffff8431ffffdf85;
    assign coff[1132] = 64'hffff8703ffffd639;
    assign coff[1133] = 64'hffff8ce8ffffc7fd;
    assign coff[1134] = 64'hffffa035ffffab1a;
    assign coff[1135] = 64'hffff803bfffff84c;
    assign coff[1136] = 64'hffff807cfffff4df;
    assign coff[1137] = 64'hffff9df7ffffadb4;
    assign coff[1138] = 64'hffff8e73ffffc4ec;
    assign coff[1139] = 64'hffff85efffffd97c;
    assign coff[1140] = 64'hffff851bffffdc35;
    assign coff[1141] = 64'hffff8fcbffffc269;
    assign coff[1142] = 64'hffff9c28ffffafe7;
    assign coff[1143] = 64'hffff80c4fffff20a;
    assign coff[1144] = 64'hffff8231ffffe86d;
    assign coff[1145] = 64'hffff965fffffb7b5;
    assign coff[1146] = 64'hffff94caffffba13;
    assign coff[1147] = 64'hffff82bfffffe5a2;
    assign coff[1148] = 64'hffff8935ffffd056;
    assign coff[1149] = 64'hffff8a4cffffcdb4;
    assign coff[1150] = 64'hffffa47dffffa681;
    assign coff[1151] = 64'hffff8002fffffe94;
    assign coff[1152] = 64'hffff8001ffffff11;
    assign coff[1153] = 64'hffffa4d5ffffa627;
    assign coff[1154] = 64'hffff8a1affffce28;
    assign coff[1155] = 64'hffff8964ffffcfe1;
    assign coff[1156] = 64'hffff82a5ffffe61d;
    assign coff[1157] = 64'hffff950effffb9aa;
    assign coff[1158] = 64'hffff9618ffffb81d;
    assign coff[1159] = 64'hffff8248ffffe7f2;
    assign coff[1160] = 64'hffff80b6fffff287;
    assign coff[1161] = 64'hffff9c77ffffaf85;
    assign coff[1162] = 64'hffff8f8fffffc2d7;
    assign coff[1163] = 64'hffff853fffffdbbd;
    assign coff[1164] = 64'hffff85c9ffffd9f4;
    assign coff[1165] = 64'hffff8eadffffc47c;
    assign coff[1166] = 64'hffff9da6ffffae14;
    assign coff[1167] = 64'hffff8087fffff462;
    assign coff[1168] = 64'hffff8034fffff8ca;
    assign coff[1169] = 64'hffffa089ffffaabc;
    assign coff[1170] = 64'hffff8cb1ffffc86e;
    assign coff[1171] = 64'hffff872cffffd5c2;
    assign coff[1172] = 64'hffff8411ffffdfff;
    assign coff[1173] = 64'hffff91bcffffbeff;
    assign coff[1174] = 64'hffff99bfffffb301;
    assign coff[1175] = 64'hffff8140ffffee24;
    assign coff[1176] = 64'hffff8187ffffec4c;
    assign coff[1177] = 64'hffff98a3ffffb480;
    assign coff[1178] = 64'hffff92b1ffffbd66;
    assign coff[1179] = 64'hffff839dffffe1ce;
    assign coff[1180] = 64'hffff87cdffffd400;
    assign coff[1181] = 64'hffff8be5ffffca1e;
    assign coff[1182] = 64'hffffa1c9ffffa95a;
    assign coff[1183] = 64'hffff801dfffffaa7;
    assign coff[1184] = 64'hffff8011fffffbed;
    assign coff[1185] = 64'hffffa2a8ffffa86b;
    assign coff[1186] = 64'hffff8b5dffffcb47;
    assign coff[1187] = 64'hffff883fffffd2ce;
    assign coff[1188] = 64'hffff8351ffffe30c;
    assign coff[1189] = 64'hffff935dffffbc4f;
    assign coff[1190] = 64'hffff97e4ffffb589;
    assign coff[1191] = 64'hffff81baffffeb09;
    assign coff[1192] = 64'hffff8115ffffef68;
    assign coff[1193] = 64'hffff9a85ffffb1fd;
    assign coff[1194] = 64'hffff9117ffffc019;
    assign coff[1195] = 64'hffff8464ffffdec3;
    assign coff[1196] = 64'hffff86c2ffffd6f7;
    assign coff[1197] = 64'hffff8d40ffffc749;
    assign coff[1198] = 64'hffff9fb0ffffabb1;
    assign coff[1199] = 64'hffff8048fffff784;
    assign coff[1200] = 64'hffff806bfffff5a7;
    assign coff[1201] = 64'hffff9e78ffffad1a;
    assign coff[1202] = 64'hffff8e17ffffc59e;
    assign coff[1203] = 64'hffff862cffffd8bc;
    assign coff[1204] = 64'hffff84e4ffffdcf6;
    assign coff[1205] = 64'hffff902cffffc1b9;
    assign coff[1206] = 64'hffff9babffffb084;
    assign coff[1207] = 64'hffff80dafffff142;
    assign coff[1208] = 64'hffff820cffffe933;
    assign coff[1209] = 64'hffff96d1ffffb710;
    assign coff[1210] = 64'hffff945cffffbabc;
    assign coff[1211] = 64'hffff82e9ffffe4de;
    assign coff[1212] = 64'hffff88eaffffd111;
    assign coff[1213] = 64'hffff8a9bffffccfc;
    assign coff[1214] = 64'hffffa3f1ffffa711;
    assign coff[1215] = 64'hffff8005fffffdcb;
    assign coff[1216] = 64'hffff8006fffffd7f;
    assign coff[1217] = 64'hffffa3bdffffa747;
    assign coff[1218] = 64'hffff8ab9ffffccb7;
    assign coff[1219] = 64'hffff88cfffffd157;
    assign coff[1220] = 64'hffff82f9ffffe494;
    assign coff[1221] = 64'hffff9434ffffbafb;
    assign coff[1222] = 64'hffff96fcffffb6d2;
    assign coff[1223] = 64'hffff81ffffffe97d;
    assign coff[1224] = 64'hffff80e3fffff0f7;
    assign coff[1225] = 64'hffff9b7cffffb0c0;
    assign coff[1226] = 64'hffff9051ffffc177;
    assign coff[1227] = 64'hffff84cfffffdd3f;
    assign coff[1228] = 64'hffff8643ffffd875;
    assign coff[1229] = 64'hffff8df5ffffc5e1;
    assign coff[1230] = 64'hffff9ea9fffface1;
    assign coff[1231] = 64'hffff8065fffff5f3;
    assign coff[1232] = 64'hffff804dfffff738;
    assign coff[1233] = 64'hffff9f7fffffabe9;
    assign coff[1234] = 64'hffff8d62ffffc705;
    assign coff[1235] = 64'hffff86a9ffffd73e;
    assign coff[1236] = 64'hffff8478ffffde7a;
    assign coff[1237] = 64'hffff90f2ffffc05b;
    assign coff[1238] = 64'hffff9ab3ffffb1c1;
    assign coff[1239] = 64'hffff810bffffefb3;
    assign coff[1240] = 64'hffff81c7ffffeabf;
    assign coff[1241] = 64'hffff97b8ffffb5c7;
    assign coff[1242] = 64'hffff9385ffffbc0f;
    assign coff[1243] = 64'hffff8340ffffe355;
    assign coff[1244] = 64'hffff8859ffffd288;
    assign coff[1245] = 64'hffff8b3effffcb8c;
    assign coff[1246] = 64'hffffa2dcffffa834;
    assign coff[1247] = 64'hffff800efffffc39;
    assign coff[1248] = 64'hffff8020fffffa5b;
    assign coff[1249] = 64'hffffa197ffffa992;
    assign coff[1250] = 64'hffff8c05ffffc9da;
    assign coff[1251] = 64'hffff87b3ffffd447;
    assign coff[1252] = 64'hffff83afffffe185;
    assign coff[1253] = 64'hffff928affffbda6;
    assign coff[1254] = 64'hffff98d0ffffb444;
    assign coff[1255] = 64'hffff817bffffec96;
    assign coff[1256] = 64'hffff814bffffedda;
    assign coff[1257] = 64'hffff9992ffffb33d;
    assign coff[1258] = 64'hffff91e2ffffbebe;
    assign coff[1259] = 64'hffff83feffffe048;
    assign coff[1260] = 64'hffff8745ffffd57b;
    assign coff[1261] = 64'hffff8c90ffffc8b2;
    assign coff[1262] = 64'hffffa0bbffffaa84;
    assign coff[1263] = 64'hffff8030fffff915;
    assign coff[1264] = 64'hffff808efffff417;
    assign coff[1265] = 64'hffff9d76ffffae4e;
    assign coff[1266] = 64'hffff8ed1ffffc43a;
    assign coff[1267] = 64'hffff85b3ffffda3c;
    assign coff[1268] = 64'hffff8554ffffdb74;
    assign coff[1269] = 64'hffff8f6bffffc319;
    assign coff[1270] = 64'hffff9ca7ffffaf4b;
    assign coff[1271] = 64'hffff80aefffff2d2;
    assign coff[1272] = 64'hffff8256ffffe7a8;
    assign coff[1273] = 64'hffff95eeffffb85b;
    assign coff[1274] = 64'hffff9538ffffb96b;
    assign coff[1275] = 64'hffff8296ffffe667;
    assign coff[1276] = 64'hffff8980ffffcf9b;
    assign coff[1277] = 64'hffff89fdffffce6d;
    assign coff[1278] = 64'hffffa50affffa5f1;
    assign coff[1279] = 64'hffff8000ffffff5d;
    assign coff[1280] = 64'hffff8000ffffff76;
    assign coff[1281] = 64'hffffa51cffffa5df;
    assign coff[1282] = 64'hffff89f3ffffce85;
    assign coff[1283] = 64'hffff898affffcf84;
    assign coff[1284] = 64'hffff8291ffffe680;
    assign coff[1285] = 64'hffff9546ffffb956;
    assign coff[1286] = 64'hffff95dfffffb870;
    assign coff[1287] = 64'hffff825bffffe78f;
    assign coff[1288] = 64'hffff80acfffff2eb;
    assign coff[1289] = 64'hffff9cb7ffffaf37;
    assign coff[1290] = 64'hffff8f5fffffc330;
    assign coff[1291] = 64'hffff855bffffdb5c;
    assign coff[1292] = 64'hffff85abffffda54;
    assign coff[1293] = 64'hffff8edcffffc423;
    assign coff[1294] = 64'hffff9d66ffffae62;
    assign coff[1295] = 64'hffff8091fffff3fe;
    assign coff[1296] = 64'hffff802ffffff92e;
    assign coff[1297] = 64'hffffa0ccffffaa71;
    assign coff[1298] = 64'hffff8c85ffffc8c9;
    assign coff[1299] = 64'hffff874dffffd563;
    assign coff[1300] = 64'hffff83f8ffffe060;
    assign coff[1301] = 64'hffff91efffffbea9;
    assign coff[1302] = 64'hffff9983ffffb351;
    assign coff[1303] = 64'hffff814fffffedc1;
    assign coff[1304] = 64'hffff8177ffffecaf;
    assign coff[1305] = 64'hffff98deffffb42f;
    assign coff[1306] = 64'hffff927dffffbdbb;
    assign coff[1307] = 64'hffff83b5ffffe16c;
    assign coff[1308] = 64'hffff87aaffffd45f;
    assign coff[1309] = 64'hffff8c0fffffc9c3;
    assign coff[1310] = 64'hffffa186ffffa9a4;
    assign coff[1311] = 64'hffff8021fffffa42;
    assign coff[1312] = 64'hffff800efffffc52;
    assign coff[1313] = 64'hffffa2edffffa821;
    assign coff[1314] = 64'hffff8b33ffffcba3;
    assign coff[1315] = 64'hffff8862ffffd270;
    assign coff[1316] = 64'hffff833bffffe36e;
    assign coff[1317] = 64'hffff9392ffffbbfa;
    assign coff[1318] = 64'hffff97a9ffffb5db;
    assign coff[1319] = 64'hffff81cbffffeaa6;
    assign coff[1320] = 64'hffff8108ffffefcc;
    assign coff[1321] = 64'hffff9ac3ffffb1ad;
    assign coff[1322] = 64'hffff90e5ffffc071;
    assign coff[1323] = 64'hffff847effffde62;
    assign coff[1324] = 64'hffff86a1ffffd756;
    assign coff[1325] = 64'hffff8d6dffffc6ef;
    assign coff[1326] = 64'hffff9f6effffabfc;
    assign coff[1327] = 64'hffff804ffffff71f;
    assign coff[1328] = 64'hffff8063fffff60c;
    assign coff[1329] = 64'hffff9ebaffffacce;
    assign coff[1330] = 64'hffff8de9ffffc5f8;
    assign coff[1331] = 64'hffff864bffffd85d;
    assign coff[1332] = 64'hffff84c8ffffdd57;
    assign coff[1333] = 64'hffff905dffffc161;
    assign coff[1334] = 64'hffff9b6dffffb0d3;
    assign coff[1335] = 64'hffff80e6fffff0de;
    assign coff[1336] = 64'hffff81faffffe996;
    assign coff[1337] = 64'hffff970affffb6bd;
    assign coff[1338] = 64'hffff9426ffffbb11;
    assign coff[1339] = 64'hffff82feffffe47b;
    assign coff[1340] = 64'hffff88c6ffffd16e;
    assign coff[1341] = 64'hffff8ac3ffffcca0;
    assign coff[1342] = 64'hffffa3abffffa759;
    assign coff[1343] = 64'hffff8007fffffd66;
    assign coff[1344] = 64'hffff8004fffffde4;
    assign coff[1345] = 64'hffffa403ffffa6ff;
    assign coff[1346] = 64'hffff8a91ffffcd13;
    assign coff[1347] = 64'hffff88f4ffffd0f9;
    assign coff[1348] = 64'hffff82e3ffffe4f6;
    assign coff[1349] = 64'hffff946affffbaa7;
    assign coff[1350] = 64'hffff96c2ffffb724;
    assign coff[1351] = 64'hffff8211ffffe91a;
    assign coff[1352] = 64'hffff80d7fffff15b;
    assign coff[1353] = 64'hffff9bbbffffb071;
    assign coff[1354] = 64'hffff9020ffffc1cf;
    assign coff[1355] = 64'hffff84eaffffdcde;
    assign coff[1356] = 64'hffff8624ffffd8d4;
    assign coff[1357] = 64'hffff8e22ffffc588;
    assign coff[1358] = 64'hffff9e68ffffad2d;
    assign coff[1359] = 64'hffff806dfffff58e;
    assign coff[1360] = 64'hffff8046fffff79d;
    assign coff[1361] = 64'hffff9fc1ffffab9e;
    assign coff[1362] = 64'hffff8d35ffffc75f;
    assign coff[1363] = 64'hffff86caffffd6df;
    assign coff[1364] = 64'hffff845effffdedb;
    assign coff[1365] = 64'hffff9124ffffc004;
    assign coff[1366] = 64'hffff9a76ffffb211;
    assign coff[1367] = 64'hffff8118ffffef4f;
    assign coff[1368] = 64'hffff81b6ffffeb22;
    assign coff[1369] = 64'hffff97f2ffffb575;
    assign coff[1370] = 64'hffff9350ffffbc65;
    assign coff[1371] = 64'hffff8357ffffe2f3;
    assign coff[1372] = 64'hffff8836ffffd2e6;
    assign coff[1373] = 64'hffff8b67ffffcb30;
    assign coff[1374] = 64'hffffa297ffffa87d;
    assign coff[1375] = 64'hffff8011fffffbd4;
    assign coff[1376] = 64'hffff801cfffffac0;
    assign coff[1377] = 64'hffffa1dbffffa948;
    assign coff[1378] = 64'hffff8bdaffffca35;
    assign coff[1379] = 64'hffff87d5ffffd3e9;
    assign coff[1380] = 64'hffff8397ffffe1e6;
    assign coff[1381] = 64'hffff92bfffffbd50;
    assign coff[1382] = 64'hffff9894ffffb495;
    assign coff[1383] = 64'hffff818affffec33;
    assign coff[1384] = 64'hffff813dffffee3d;
    assign coff[1385] = 64'hffff99cfffffb2ed;
    assign coff[1386] = 64'hffff91afffffbf15;
    assign coff[1387] = 64'hffff8417ffffdfe6;
    assign coff[1388] = 64'hffff8724ffffd5da;
    assign coff[1389] = 64'hffff8cbcffffc858;
    assign coff[1390] = 64'hffffa078ffffaacf;
    assign coff[1391] = 64'hffff8035fffff8b1;
    assign coff[1392] = 64'hffff8085fffff47b;
    assign coff[1393] = 64'hffff9db6ffffae01;
    assign coff[1394] = 64'hffff8ea2ffffc493;
    assign coff[1395] = 64'hffff85d1ffffd9dc;
    assign coff[1396] = 64'hffff8537ffffdbd5;
    assign coff[1397] = 64'hffff8f9bffffc2c1;
    assign coff[1398] = 64'hffff9c67ffffaf99;
    assign coff[1399] = 64'hffff80b9fffff26e;
    assign coff[1400] = 64'hffff8243ffffe80a;
    assign coff[1401] = 64'hffff9626ffffb808;
    assign coff[1402] = 64'hffff9501ffffb9bf;
    assign coff[1403] = 64'hffff82aaffffe605;
    assign coff[1404] = 64'hffff895affffcff8;
    assign coff[1405] = 64'hffff8a24ffffce11;
    assign coff[1406] = 64'hffffa4c4ffffa639;
    assign coff[1407] = 64'hffff8001fffffef8;
    assign coff[1408] = 64'hffff8002fffffead;
    assign coff[1409] = 64'hffffa48fffffa66f;
    assign coff[1410] = 64'hffff8a42ffffcdcb;
    assign coff[1411] = 64'hffff893effffd03e;
    assign coff[1412] = 64'hffff82baffffe5bb;
    assign coff[1413] = 64'hffff94d7ffffb9fe;
    assign coff[1414] = 64'hffff9650ffffb7ca;
    assign coff[1415] = 64'hffff8235ffffe854;
    assign coff[1416] = 64'hffff80c1fffff223;
    assign coff[1417] = 64'hffff9c38ffffafd4;
    assign coff[1418] = 64'hffff8fbfffffc27f;
    assign coff[1419] = 64'hffff8522ffffdc1d;
    assign coff[1420] = 64'hffff85e7ffffd994;
    assign coff[1421] = 64'hffff8e7fffffc4d5;
    assign coff[1422] = 64'hffff9de7ffffadc7;
    assign coff[1423] = 64'hffff807efffff4c6;
    assign coff[1424] = 64'hffff803afffff865;
    assign coff[1425] = 64'hffffa046ffffab07;
    assign coff[1426] = 64'hffff8cddffffc814;
    assign coff[1427] = 64'hffff870bffffd621;
    assign coff[1428] = 64'hffff842affffdf9d;
    assign coff[1429] = 64'hffff9189ffffbf56;
    assign coff[1430] = 64'hffff99fcffffb2b1;
    assign coff[1431] = 64'hffff8133ffffee88;
    assign coff[1432] = 64'hffff8196ffffebe9;
    assign coff[1433] = 64'hffff9868ffffb4d2;
    assign coff[1434] = 64'hffff92e6ffffbd10;
    assign coff[1435] = 64'hffff8385ffffe230;
    assign coff[1436] = 64'hffff87efffffd3a2;
    assign coff[1437] = 64'hffff8bbbffffca79;
    assign coff[1438] = 64'hffffa20effffa910;
    assign coff[1439] = 64'hffff8019fffffb0b;
    assign coff[1440] = 64'hffff8014fffffb89;
    assign coff[1441] = 64'hffffa263ffffa8b4;
    assign coff[1442] = 64'hffff8b86ffffcaec;
    assign coff[1443] = 64'hffff881bffffd32c;
    assign coff[1444] = 64'hffff8368ffffe2aa;
    assign coff[1445] = 64'hffff9328ffffbca5;
    assign coff[1446] = 64'hffff981effffb538;
    assign coff[1447] = 64'hffff81aaffffeb6d;
    assign coff[1448] = 64'hffff8122ffffef04;
    assign coff[1449] = 64'hffff9a48ffffb24d;
    assign coff[1450] = 64'hffff914affffbfc2;
    assign coff[1451] = 64'hffff844affffdf24;
    assign coff[1452] = 64'hffff86e2ffffd698;
    assign coff[1453] = 64'hffff8d14ffffc7a3;
    assign coff[1454] = 64'hffff9ff3ffffab65;
    assign coff[1455] = 64'hffff8042fffff7e8;
    assign coff[1456] = 64'hffff8073fffff543;
    assign coff[1457] = 64'hffff9e37ffffad67;
    assign coff[1458] = 64'hffff8e45ffffc545;
    assign coff[1459] = 64'hffff860dffffd91c;
    assign coff[1460] = 64'hffff84ffffffdc96;
    assign coff[1461] = 64'hffff8ffbffffc211;
    assign coff[1462] = 64'hffff9beaffffb036;
    assign coff[1463] = 64'hffff80cffffff1a6;
    assign coff[1464] = 64'hffff821effffe8d0;
    assign coff[1465] = 64'hffff9697ffffb762;
    assign coff[1466] = 64'hffff9493ffffba67;
    assign coff[1467] = 64'hffff82d4ffffe540;
    assign coff[1468] = 64'hffff890fffffd0b3;
    assign coff[1469] = 64'hffff8a73ffffcd58;
    assign coff[1470] = 64'hffffa437ffffa6c9;
    assign coff[1471] = 64'hffff8003fffffe2f;
    assign coff[1472] = 64'hffff8008fffffd1b;
    assign coff[1473] = 64'hffffa377ffffa790;
    assign coff[1474] = 64'hffff8ae2ffffcc5b;
    assign coff[1475] = 64'hffff88aaffffd1b4;
    assign coff[1476] = 64'hffff830effffe432;
    assign coff[1477] = 64'hffff93feffffbb50;
    assign coff[1478] = 64'hffff9735ffffb67f;
    assign coff[1479] = 64'hffff81edffffe9e0;
    assign coff[1480] = 64'hffff80effffff093;
    assign coff[1481] = 64'hffff9b3effffb10f;
    assign coff[1482] = 64'hffff9082ffffc11f;
    assign coff[1483] = 64'hffff84b4ffffdda0;
    assign coff[1484] = 64'hffff8662ffffd815;
    assign coff[1485] = 64'hffff8dc7ffffc63b;
    assign coff[1486] = 64'hffff9eebffffac94;
    assign coff[1487] = 64'hffff805dfffff657;
    assign coff[1488] = 64'hffff8054fffff6d4;
    assign coff[1489] = 64'hffff9f3dffffac35;
    assign coff[1490] = 64'hffff8d8fffffc6ab;
    assign coff[1491] = 64'hffff868affffd79e;
    assign coff[1492] = 64'hffff8492ffffde19;
    assign coff[1493] = 64'hffff90c0ffffc0b2;
    assign coff[1494] = 64'hffff9af1ffffb172;
    assign coff[1495] = 64'hffff80fefffff016;
    assign coff[1496] = 64'hffff81d8ffffea5c;
    assign coff[1497] = 64'hffff977effffb619;
    assign coff[1498] = 64'hffff93baffffbbba;
    assign coff[1499] = 64'hffff832affffe3b7;
    assign coff[1500] = 64'hffff887dffffd22a;
    assign coff[1501] = 64'hffff8b15ffffcbe8;
    assign coff[1502] = 64'hffffa321ffffa7eb;
    assign coff[1503] = 64'hffff800bfffffc9d;
    assign coff[1504] = 64'hffff8024fffff9f7;
    assign coff[1505] = 64'hffffa153ffffa9dc;
    assign coff[1506] = 64'hffff8c2fffffc97f;
    assign coff[1507] = 64'hffff8791ffffd4a6;
    assign coff[1508] = 64'hffff83c7ffffe123;
    assign coff[1509] = 64'hffff9256ffffbdfc;
    assign coff[1510] = 64'hffff990bffffb3f3;
    assign coff[1511] = 64'hffff816cffffecfa;
    assign coff[1512] = 64'hffff815affffed76;
    assign coff[1513] = 64'hffff9956ffffb38e;
    assign coff[1514] = 64'hffff9216ffffbe68;
    assign coff[1515] = 64'hffff83e5ffffe0a9;
    assign coff[1516] = 64'hffff8766ffffd51c;
    assign coff[1517] = 64'hffff8c65ffffc90d;
    assign coff[1518] = 64'hffffa0feffffaa39;
    assign coff[1519] = 64'hffff802bfffff979;
    assign coff[1520] = 64'hffff8098fffff3b3;
    assign coff[1521] = 64'hffff9d36ffffae9c;
    assign coff[1522] = 64'hffff8f00ffffc3e1;
    assign coff[1523] = 64'hffff8595ffffda9c;
    assign coff[1524] = 64'hffff8571ffffdb14;
    assign coff[1525] = 64'hffff8f3bffffc372;
    assign coff[1526] = 64'hffff9ce6ffffaefd;
    assign coff[1527] = 64'hffff80a4fffff336;
    assign coff[1528] = 64'hffff8269ffffe745;
    assign coff[1529] = 64'hffff95b5ffffb8af;
    assign coff[1530] = 64'hffff9570ffffb917;
    assign coff[1531] = 64'hffff8282ffffe6ca;
    assign coff[1532] = 64'hffff89a6ffffcf3e;
    assign coff[1533] = 64'hffff89d6ffffceca;
    assign coff[1534] = 64'hffffa551ffffa5aa;
    assign coff[1535] = 64'hffff8000ffffffc1;
    assign coff[1536] = 64'hffff8000ffffffa8;
    assign coff[1537] = 64'hffffa53fffffa5bc;
    assign coff[1538] = 64'hffff89e0ffffceb3;
    assign coff[1539] = 64'hffff899dffffcf56;
    assign coff[1540] = 64'hffff8287ffffe6b1;
    assign coff[1541] = 64'hffff9562ffffb92c;
    assign coff[1542] = 64'hffff95c3ffffb89a;
    assign coff[1543] = 64'hffff8265ffffe75e;
    assign coff[1544] = 64'hffff80a7fffff31d;
    assign coff[1545] = 64'hffff9cd6ffffaf10;
    assign coff[1546] = 64'hffff8f47ffffc35c;
    assign coff[1547] = 64'hffff856affffdb2c;
    assign coff[1548] = 64'hffff859dffffda84;
    assign coff[1549] = 64'hffff8ef4ffffc3f7;
    assign coff[1550] = 64'hffff9d46ffffae88;
    assign coff[1551] = 64'hffff8095fffff3cc;
    assign coff[1552] = 64'hffff802cfffff960;
    assign coff[1553] = 64'hffffa0eeffffaa4c;
    assign coff[1554] = 64'hffff8c70ffffc8f6;
    assign coff[1555] = 64'hffff875effffd534;
    assign coff[1556] = 64'hffff83ecffffe091;
    assign coff[1557] = 64'hffff9209ffffbe7d;
    assign coff[1558] = 64'hffff9965ffffb37a;
    assign coff[1559] = 64'hffff8156ffffed8f;
    assign coff[1560] = 64'hffff8170ffffece1;
    assign coff[1561] = 64'hffff98fcffffb407;
    assign coff[1562] = 64'hffff9263ffffbde6;
    assign coff[1563] = 64'hffff83c1ffffe13b;
    assign coff[1564] = 64'hffff8799ffffd48e;
    assign coff[1565] = 64'hffff8c25ffffc995;
    assign coff[1566] = 64'hffffa164ffffa9c9;
    assign coff[1567] = 64'hffff8023fffffa10;
    assign coff[1568] = 64'hffff800cfffffc84;
    assign coff[1569] = 64'hffffa30fffffa7fd;
    assign coff[1570] = 64'hffff8b1fffffcbd1;
    assign coff[1571] = 64'hffff8874ffffd241;
    assign coff[1572] = 64'hffff8330ffffe39f;
    assign coff[1573] = 64'hffff93adffffbbd0;
    assign coff[1574] = 64'hffff978cffffb604;
    assign coff[1575] = 64'hffff81d3ffffea75;
    assign coff[1576] = 64'hffff8101ffffeffe;
    assign coff[1577] = 64'hffff9ae1ffffb186;
    assign coff[1578] = 64'hffff90ccffffc09c;
    assign coff[1579] = 64'hffff848cffffde31;
    assign coff[1580] = 64'hffff8692ffffd786;
    assign coff[1581] = 64'hffff8d83ffffc6c2;
    assign coff[1582] = 64'hffff9f4dffffac22;
    assign coff[1583] = 64'hffff8052fffff6ed;
    assign coff[1584] = 64'hffff805ffffff63e;
    assign coff[1585] = 64'hffff9edaffffaca8;
    assign coff[1586] = 64'hffff8dd2ffffc625;
    assign coff[1587] = 64'hffff865affffd82d;
    assign coff[1588] = 64'hffff84bbffffdd88;
    assign coff[1589] = 64'hffff9076ffffc135;
    assign coff[1590] = 64'hffff9b4effffb0fb;
    assign coff[1591] = 64'hffff80ecfffff0ac;
    assign coff[1592] = 64'hffff81f2ffffe9c7;
    assign coff[1593] = 64'hffff9727ffffb694;
    assign coff[1594] = 64'hffff940bffffbb3b;
    assign coff[1595] = 64'hffff8309ffffe44a;
    assign coff[1596] = 64'hffff88b3ffffd19d;
    assign coff[1597] = 64'hffff8ad8ffffcc72;
    assign coff[1598] = 64'hffffa389ffffa77e;
    assign coff[1599] = 64'hffff8008fffffd34;
    assign coff[1600] = 64'hffff8004fffffe16;
    assign coff[1601] = 64'hffffa426ffffa6db;
    assign coff[1602] = 64'hffff8a7dffffcd41;
    assign coff[1603] = 64'hffff8906ffffd0ca;
    assign coff[1604] = 64'hffff82d9ffffe527;
    assign coff[1605] = 64'hffff9485ffffba7d;
    assign coff[1606] = 64'hffff96a6ffffb74e;
    assign coff[1607] = 64'hffff821affffe8e9;
    assign coff[1608] = 64'hffff80d1fffff18d;
    assign coff[1609] = 64'hffff9bdaffffb049;
    assign coff[1610] = 64'hffff9007ffffc1fb;
    assign coff[1611] = 64'hffff84f8ffffdcae;
    assign coff[1612] = 64'hffff8615ffffd904;
    assign coff[1613] = 64'hffff8e39ffffc55b;
    assign coff[1614] = 64'hffff9e48ffffad54;
    assign coff[1615] = 64'hffff8071fffff55c;
    assign coff[1616] = 64'hffff8043fffff7cf;
    assign coff[1617] = 64'hffff9fe2ffffab78;
    assign coff[1618] = 64'hffff8d1fffffc78c;
    assign coff[1619] = 64'hffff86daffffd6af;
    assign coff[1620] = 64'hffff8451ffffdf0c;
    assign coff[1621] = 64'hffff913dffffbfd8;
    assign coff[1622] = 64'hffff9a57ffffb239;
    assign coff[1623] = 64'hffff811effffef1d;
    assign coff[1624] = 64'hffff81aeffffeb54;
    assign coff[1625] = 64'hffff9810ffffb54c;
    assign coff[1626] = 64'hffff9335ffffbc8f;
    assign coff[1627] = 64'hffff8362ffffe2c2;
    assign coff[1628] = 64'hffff8824ffffd315;
    assign coff[1629] = 64'hffff8b7cffffcb02;
    assign coff[1630] = 64'hffffa274ffffa8a2;
    assign coff[1631] = 64'hffff8013fffffba2;
    assign coff[1632] = 64'hffff801afffffaf2;
    assign coff[1633] = 64'hffffa1fdffffa923;
    assign coff[1634] = 64'hffff8bc5ffffca63;
    assign coff[1635] = 64'hffff87e7ffffd3ba;
    assign coff[1636] = 64'hffff838bffffe217;
    assign coff[1637] = 64'hffff92d9ffffbd25;
    assign coff[1638] = 64'hffff9877ffffb4bd;
    assign coff[1639] = 64'hffff8192ffffec01;
    assign coff[1640] = 64'hffff8136ffffee6f;
    assign coff[1641] = 64'hffff99edffffb2c5;
    assign coff[1642] = 64'hffff9196ffffbf40;
    assign coff[1643] = 64'hffff8424ffffdfb6;
    assign coff[1644] = 64'hffff8713ffffd609;
    assign coff[1645] = 64'hffff8cd2ffffc82b;
    assign coff[1646] = 64'hffffa057ffffaaf4;
    assign coff[1647] = 64'hffff8038fffff87e;
    assign coff[1648] = 64'hffff8080fffff4ad;
    assign coff[1649] = 64'hffff9dd6ffffadda;
    assign coff[1650] = 64'hffff8e8affffc4bf;
    assign coff[1651] = 64'hffff85e0ffffd9ac;
    assign coff[1652] = 64'hffff8529ffffdc05;
    assign coff[1653] = 64'hffff8fb3ffffc295;
    assign coff[1654] = 64'hffff9c48ffffafc0;
    assign coff[1655] = 64'hffff80befffff23c;
    assign coff[1656] = 64'hffff823affffe83c;
    assign coff[1657] = 64'hffff9642ffffb7df;
    assign coff[1658] = 64'hffff94e5ffffb9e9;
    assign coff[1659] = 64'hffff82b4ffffe5d3;
    assign coff[1660] = 64'hffff8947ffffd027;
    assign coff[1661] = 64'hffff8a38ffffcde3;
    assign coff[1662] = 64'hffffa4a0ffffa65d;
    assign coff[1663] = 64'hffff8002fffffec6;
    assign coff[1664] = 64'hffff8001fffffedf;
    assign coff[1665] = 64'hffffa4b2ffffa64b;
    assign coff[1666] = 64'hffff8a2effffcdfa;
    assign coff[1667] = 64'hffff8951ffffd010;
    assign coff[1668] = 64'hffff82afffffe5ec;
    assign coff[1669] = 64'hffff94f3ffffb9d4;
    assign coff[1670] = 64'hffff9634ffffb7f3;
    assign coff[1671] = 64'hffff823effffe823;
    assign coff[1672] = 64'hffff80bbfffff255;
    assign coff[1673] = 64'hffff9c58ffffafac;
    assign coff[1674] = 64'hffff8fa7ffffc2ab;
    assign coff[1675] = 64'hffff8530ffffdbed;
    assign coff[1676] = 64'hffff85d8ffffd9c4;
    assign coff[1677] = 64'hffff8e96ffffc4a9;
    assign coff[1678] = 64'hffff9dc6ffffadee;
    assign coff[1679] = 64'hffff8083fffff494;
    assign coff[1680] = 64'hffff8037fffff898;
    assign coff[1681] = 64'hffffa067ffffaae1;
    assign coff[1682] = 64'hffff8cc7ffffc841;
    assign coff[1683] = 64'hffff871bffffd5f1;
    assign coff[1684] = 64'hffff841dffffdfce;
    assign coff[1685] = 64'hffff91a2ffffbf2a;
    assign coff[1686] = 64'hffff99deffffb2d9;
    assign coff[1687] = 64'hffff813affffee56;
    assign coff[1688] = 64'hffff818effffec1a;
    assign coff[1689] = 64'hffff9885ffffb4a9;
    assign coff[1690] = 64'hffff92ccffffbd3b;
    assign coff[1691] = 64'hffff8391ffffe1ff;
    assign coff[1692] = 64'hffff87deffffd3d1;
    assign coff[1693] = 64'hffff8bd0ffffca4c;
    assign coff[1694] = 64'hffffa1ecffffa935;
    assign coff[1695] = 64'hffff801bfffffad9;
    assign coff[1696] = 64'hffff8012fffffbbb;
    assign coff[1697] = 64'hffffa286ffffa88f;
    assign coff[1698] = 64'hffff8b71ffffcb19;
    assign coff[1699] = 64'hffff882dffffd2fd;
    assign coff[1700] = 64'hffff835dffffe2db;
    assign coff[1701] = 64'hffff9342ffffbc7a;
    assign coff[1702] = 64'hffff9801ffffb560;
    assign coff[1703] = 64'hffff81b2ffffeb3b;
    assign coff[1704] = 64'hffff811bffffef36;
    assign coff[1705] = 64'hffff9a67ffffb225;
    assign coff[1706] = 64'hffff9131ffffbfee;
    assign coff[1707] = 64'hffff8457ffffdef3;
    assign coff[1708] = 64'hffff86d2ffffd6c7;
    assign coff[1709] = 64'hffff8d2affffc776;
    assign coff[1710] = 64'hffff9fd2ffffab8b;
    assign coff[1711] = 64'hffff8045fffff7b6;
    assign coff[1712] = 64'hffff806ffffff575;
    assign coff[1713] = 64'hffff9e58ffffad41;
    assign coff[1714] = 64'hffff8e2effffc572;
    assign coff[1715] = 64'hffff861cffffd8ec;
    assign coff[1716] = 64'hffff84f1ffffdcc6;
    assign coff[1717] = 64'hffff9014ffffc1e5;
    assign coff[1718] = 64'hffff9bcaffffb05d;
    assign coff[1719] = 64'hffff80d4fffff174;
    assign coff[1720] = 64'hffff8215ffffe901;
    assign coff[1721] = 64'hffff96b4ffffb739;
    assign coff[1722] = 64'hffff9478ffffba92;
    assign coff[1723] = 64'hffff82deffffe50f;
    assign coff[1724] = 64'hffff88fdffffd0e2;
    assign coff[1725] = 64'hffff8a87ffffcd2a;
    assign coff[1726] = 64'hffffa414ffffa6ed;
    assign coff[1727] = 64'hffff8004fffffdfd;
    assign coff[1728] = 64'hffff8007fffffd4d;
    assign coff[1729] = 64'hffffa39affffa76b;
    assign coff[1730] = 64'hffff8aceffffcc89;
    assign coff[1731] = 64'hffff88bdffffd186;
    assign coff[1732] = 64'hffff8304ffffe463;
    assign coff[1733] = 64'hffff9419ffffbb26;
    assign coff[1734] = 64'hffff9718ffffb6a8;
    assign coff[1735] = 64'hffff81f6ffffe9af;
    assign coff[1736] = 64'hffff80e9fffff0c5;
    assign coff[1737] = 64'hffff9b5dffffb0e7;
    assign coff[1738] = 64'hffff9069ffffc14b;
    assign coff[1739] = 64'hffff84c1ffffdd6f;
    assign coff[1740] = 64'hffff8653ffffd845;
    assign coff[1741] = 64'hffff8ddeffffc60e;
    assign coff[1742] = 64'hffff9ecaffffacbb;
    assign coff[1743] = 64'hffff8061fffff625;
    assign coff[1744] = 64'hffff8051fffff706;
    assign coff[1745] = 64'hffff9f5effffac0f;
    assign coff[1746] = 64'hffff8d78ffffc6d8;
    assign coff[1747] = 64'hffff869affffd76e;
    assign coff[1748] = 64'hffff8485ffffde49;
    assign coff[1749] = 64'hffff90d9ffffc086;
    assign coff[1750] = 64'hffff9ad2ffffb199;
    assign coff[1751] = 64'hffff8104ffffefe5;
    assign coff[1752] = 64'hffff81cfffffea8d;
    assign coff[1753] = 64'hffff979bffffb5f0;
    assign coff[1754] = 64'hffff939fffffbbe5;
    assign coff[1755] = 64'hffff8335ffffe386;
    assign coff[1756] = 64'hffff886bffffd259;
    assign coff[1757] = 64'hffff8b29ffffcbba;
    assign coff[1758] = 64'hffffa2feffffa80f;
    assign coff[1759] = 64'hffff800dfffffc6b;
    assign coff[1760] = 64'hffff8022fffffa29;
    assign coff[1761] = 64'hffffa175ffffa9b7;
    assign coff[1762] = 64'hffff8c1affffc9ac;
    assign coff[1763] = 64'hffff87a2ffffd476;
    assign coff[1764] = 64'hffff83bbffffe154;
    assign coff[1765] = 64'hffff9270ffffbdd1;
    assign coff[1766] = 64'hffff98edffffb41b;
    assign coff[1767] = 64'hffff8173ffffecc8;
    assign coff[1768] = 64'hffff8152ffffeda8;
    assign coff[1769] = 64'hffff9974ffffb365;
    assign coff[1770] = 64'hffff91fcffffbe93;
    assign coff[1771] = 64'hffff83f2ffffe078;
    assign coff[1772] = 64'hffff8756ffffd54b;
    assign coff[1773] = 64'hffff8c7bffffc8e0;
    assign coff[1774] = 64'hffffa0ddffffaa5e;
    assign coff[1775] = 64'hffff802dfffff947;
    assign coff[1776] = 64'hffff8093fffff3e5;
    assign coff[1777] = 64'hffff9d56ffffae75;
    assign coff[1778] = 64'hffff8ee8ffffc40d;
    assign coff[1779] = 64'hffff85a4ffffda6c;
    assign coff[1780] = 64'hffff8562ffffdb44;
    assign coff[1781] = 64'hffff8f53ffffc346;
    assign coff[1782] = 64'hffff9cc6ffffaf24;
    assign coff[1783] = 64'hffff80a9fffff304;
    assign coff[1784] = 64'hffff8260ffffe776;
    assign coff[1785] = 64'hffff95d1ffffb885;
    assign coff[1786] = 64'hffff9554ffffb941;
    assign coff[1787] = 64'hffff828cffffe698;
    assign coff[1788] = 64'hffff8993ffffcf6d;
    assign coff[1789] = 64'hffff89eaffffce9c;
    assign coff[1790] = 64'hffffa52effffa5ce;
    assign coff[1791] = 64'hffff8000ffffff8f;
    assign coff[1792] = 64'hffff8001ffffff44;
    assign coff[1793] = 64'hffffa4f9ffffa603;
    assign coff[1794] = 64'hffff8a07ffffce56;
    assign coff[1795] = 64'hffff8977ffffcfb3;
    assign coff[1796] = 64'hffff829bffffe64f;
    assign coff[1797] = 64'hffff952affffb980;
    assign coff[1798] = 64'hffff95fcffffb847;
    assign coff[1799] = 64'hffff8251ffffe7c0;
    assign coff[1800] = 64'hffff80b1fffff2b9;
    assign coff[1801] = 64'hffff9c97ffffaf5e;
    assign coff[1802] = 64'hffff8f77ffffc303;
    assign coff[1803] = 64'hffff854dffffdb8c;
    assign coff[1804] = 64'hffff85baffffda24;
    assign coff[1805] = 64'hffff8ec5ffffc450;
    assign coff[1806] = 64'hffff9d86ffffae3b;
    assign coff[1807] = 64'hffff808cfffff430;
    assign coff[1808] = 64'hffff8031fffff8fc;
    assign coff[1809] = 64'hffffa0aaffffaa96;
    assign coff[1810] = 64'hffff8c9bffffc89c;
    assign coff[1811] = 64'hffff873cffffd592;
    assign coff[1812] = 64'hffff8404ffffe02f;
    assign coff[1813] = 64'hffff91d6ffffbed4;
    assign coff[1814] = 64'hffff99a1ffffb329;
    assign coff[1815] = 64'hffff8148ffffedf2;
    assign coff[1816] = 64'hffff817fffffec7e;
    assign coff[1817] = 64'hffff98c1ffffb458;
    assign coff[1818] = 64'hffff9297ffffbd90;
    assign coff[1819] = 64'hffff83a9ffffe19d;
    assign coff[1820] = 64'hffff87bbffffd430;
    assign coff[1821] = 64'hffff8bfaffffc9f1;
    assign coff[1822] = 64'hffffa1a8ffffa97f;
    assign coff[1823] = 64'hffff801ffffffa74;
    assign coff[1824] = 64'hffff800ffffffc1f;
    assign coff[1825] = 64'hffffa2caffffa846;
    assign coff[1826] = 64'hffff8b48ffffcb75;
    assign coff[1827] = 64'hffff8850ffffd29f;
    assign coff[1828] = 64'hffff8346ffffe33d;
    assign coff[1829] = 64'hffff9377ffffbc25;
    assign coff[1830] = 64'hffff97c6ffffb5b2;
    assign coff[1831] = 64'hffff81c3ffffead8;
    assign coff[1832] = 64'hffff810effffef9a;
    assign coff[1833] = 64'hffff9aa4ffffb1d5;
    assign coff[1834] = 64'hffff90feffffc045;
    assign coff[1835] = 64'hffff8471ffffde92;
    assign coff[1836] = 64'hffff86b2ffffd726;
    assign coff[1837] = 64'hffff8d57ffffc71c;
    assign coff[1838] = 64'hffff9f8fffffabd6;
    assign coff[1839] = 64'hffff804bfffff751;
    assign coff[1840] = 64'hffff8067fffff5d9;
    assign coff[1841] = 64'hffff9e99ffffacf4;
    assign coff[1842] = 64'hffff8e00ffffc5cb;
    assign coff[1843] = 64'hffff863bffffd88c;
    assign coff[1844] = 64'hffff84d6ffffdd27;
    assign coff[1845] = 64'hffff9045ffffc18d;
    assign coff[1846] = 64'hffff9b8cffffb0ac;
    assign coff[1847] = 64'hffff80e0fffff110;
    assign coff[1848] = 64'hffff8203ffffe964;
    assign coff[1849] = 64'hffff96edffffb6e6;
    assign coff[1850] = 64'hffff9441ffffbae6;
    assign coff[1851] = 64'hffff82f3ffffe4ad;
    assign coff[1852] = 64'hffff88d8ffffd13f;
    assign coff[1853] = 64'hffff8aafffffccce;
    assign coff[1854] = 64'hffffa3ceffffa735;
    assign coff[1855] = 64'hffff8006fffffd98;
    assign coff[1856] = 64'hffff8005fffffdb1;
    assign coff[1857] = 64'hffffa3e0ffffa723;
    assign coff[1858] = 64'hffff8aa5ffffcce5;
    assign coff[1859] = 64'hffff88e1ffffd128;
    assign coff[1860] = 64'hffff82eeffffe4c5;
    assign coff[1861] = 64'hffff944fffffbad1;
    assign coff[1862] = 64'hffff96dfffffb6fb;
    assign coff[1863] = 64'hffff8208ffffe94c;
    assign coff[1864] = 64'hffff80ddfffff129;
    assign coff[1865] = 64'hffff9b9bffffb098;
    assign coff[1866] = 64'hffff9038ffffc1a3;
    assign coff[1867] = 64'hffff84ddffffdd0f;
    assign coff[1868] = 64'hffff8634ffffd8a4;
    assign coff[1869] = 64'hffff8e0bffffc5b5;
    assign coff[1870] = 64'hffff9e89ffffad07;
    assign coff[1871] = 64'hffff8069fffff5c0;
    assign coff[1872] = 64'hffff804afffff76b;
    assign coff[1873] = 64'hffff9fa0ffffabc4;
    assign coff[1874] = 64'hffff8d4bffffc732;
    assign coff[1875] = 64'hffff86baffffd70f;
    assign coff[1876] = 64'hffff846bffffdeaa;
    assign coff[1877] = 64'hffff910bffffc02f;
    assign coff[1878] = 64'hffff9a95ffffb1e9;
    assign coff[1879] = 64'hffff8111ffffef81;
    assign coff[1880] = 64'hffff81bfffffeaf1;
    assign coff[1881] = 64'hffff97d5ffffb59e;
    assign coff[1882] = 64'hffff936affffbc3a;
    assign coff[1883] = 64'hffff834cffffe324;
    assign coff[1884] = 64'hffff8847ffffd2b7;
    assign coff[1885] = 64'hffff8b52ffffcb5e;
    assign coff[1886] = 64'hffffa2b9ffffa858;
    assign coff[1887] = 64'hffff8010fffffc06;
    assign coff[1888] = 64'hffff801efffffa8e;
    assign coff[1889] = 64'hffffa1b8ffffa96d;
    assign coff[1890] = 64'hffff8befffffca07;
    assign coff[1891] = 64'hffff87c4ffffd418;
    assign coff[1892] = 64'hffff83a3ffffe1b5;
    assign coff[1893] = 64'hffff92a4ffffbd7b;
    assign coff[1894] = 64'hffff98b2ffffb46c;
    assign coff[1895] = 64'hffff8183ffffec65;
    assign coff[1896] = 64'hffff8144ffffee0b;
    assign coff[1897] = 64'hffff99b0ffffb315;
    assign coff[1898] = 64'hffff91c9ffffbee9;
    assign coff[1899] = 64'hffff840bffffe017;
    assign coff[1900] = 64'hffff8734ffffd5aa;
    assign coff[1901] = 64'hffff8ca6ffffc885;
    assign coff[1902] = 64'hffffa09affffaaa9;
    assign coff[1903] = 64'hffff8033fffff8e3;
    assign coff[1904] = 64'hffff808afffff449;
    assign coff[1905] = 64'hffff9d96ffffae28;
    assign coff[1906] = 64'hffff8eb9ffffc466;
    assign coff[1907] = 64'hffff85c2ffffda0c;
    assign coff[1908] = 64'hffff8546ffffdba5;
    assign coff[1909] = 64'hffff8f83ffffc2ed;
    assign coff[1910] = 64'hffff9c87ffffaf72;
    assign coff[1911] = 64'hffff80b3fffff2a0;
    assign coff[1912] = 64'hffff824dffffe7d9;
    assign coff[1913] = 64'hffff960affffb832;
    assign coff[1914] = 64'hffff951cffffb995;
    assign coff[1915] = 64'hffff82a0ffffe636;
    assign coff[1916] = 64'hffff896dffffcfca;
    assign coff[1917] = 64'hffff8a11ffffce3f;
    assign coff[1918] = 64'hffffa4e7ffffa615;
    assign coff[1919] = 64'hffff8001ffffff2a;
    assign coff[1920] = 64'hffff8002fffffe7a;
    assign coff[1921] = 64'hffffa46cffffa693;
    assign coff[1922] = 64'hffff8a56ffffcd9d;
    assign coff[1923] = 64'hffff892bffffd06d;
    assign coff[1924] = 64'hffff82c4ffffe58a;
    assign coff[1925] = 64'hffff94bcffffba28;
    assign coff[1926] = 64'hffff966dffffb7a0;
    assign coff[1927] = 64'hffff822cffffe886;
    assign coff[1928] = 64'hffff80c6fffff1f1;
    assign coff[1929] = 64'hffff9c19ffffaffb;
    assign coff[1930] = 64'hffff8fd7ffffc253;
    assign coff[1931] = 64'hffff8514ffffdc4d;
    assign coff[1932] = 64'hffff85f6ffffd964;
    assign coff[1933] = 64'hffff8e68ffffc502;
    assign coff[1934] = 64'hffff9e07ffffada1;
    assign coff[1935] = 64'hffff807afffff4f8;
    assign coff[1936] = 64'hffff803dfffff833;
    assign coff[1937] = 64'hffffa025ffffab2d;
    assign coff[1938] = 64'hffff8cf3ffffc7e7;
    assign coff[1939] = 64'hffff86faffffd650;
    assign coff[1940] = 64'hffff8437ffffdf6d;
    assign coff[1941] = 64'hffff9170ffffbf81;
    assign coff[1942] = 64'hffff9a1affffb289;
    assign coff[1943] = 64'hffff812cffffeeba;
    assign coff[1944] = 64'hffff819effffebb7;
    assign coff[1945] = 64'hffff984affffb4fa;
    assign coff[1946] = 64'hffff9300ffffbce5;
    assign coff[1947] = 64'hffff837affffe260;
    assign coff[1948] = 64'hffff8801ffffd373;
    assign coff[1949] = 64'hffff8ba6ffffcaa7;
    assign coff[1950] = 64'hffffa230ffffa8eb;
    assign coff[1951] = 64'hffff8017fffffb3d;
    assign coff[1952] = 64'hffff8016fffffb56;
    assign coff[1953] = 64'hffffa241ffffa8d9;
    assign coff[1954] = 64'hffff8b9bffffcabe;
    assign coff[1955] = 64'hffff880affffd35b;
    assign coff[1956] = 64'hffff8374ffffe279;
    assign coff[1957] = 64'hffff930dffffbcd0;
    assign coff[1958] = 64'hffff983cffffb50f;
    assign coff[1959] = 64'hffff81a2ffffeb9e;
    assign coff[1960] = 64'hffff8128ffffeed3;
    assign coff[1961] = 64'hffff9a2affffb275;
    assign coff[1962] = 64'hffff9163ffffbf97;
    assign coff[1963] = 64'hffff843dffffdf54;
    assign coff[1964] = 64'hffff86f2ffffd668;
    assign coff[1965] = 64'hffff8cfeffffc7d0;
    assign coff[1966] = 64'hffffa014ffffab3f;
    assign coff[1967] = 64'hffff803efffff81a;
    assign coff[1968] = 64'hffff8078fffff511;
    assign coff[1969] = 64'hffff9e17ffffad8d;
    assign coff[1970] = 64'hffff8e5cffffc518;
    assign coff[1971] = 64'hffff85feffffd94c;
    assign coff[1972] = 64'hffff850dffffdc66;
    assign coff[1973] = 64'hffff8fe3ffffc23d;
    assign coff[1974] = 64'hffff9c09ffffb00e;
    assign coff[1975] = 64'hffff80c9fffff1d8;
    assign coff[1976] = 64'hffff8227ffffe89f;
    assign coff[1977] = 64'hffff967bffffb78c;
    assign coff[1978] = 64'hffff94aeffffba3d;
    assign coff[1979] = 64'hffff82c9ffffe571;
    assign coff[1980] = 64'hffff8922ffffd084;
    assign coff[1981] = 64'hffff8a5fffffcd86;
    assign coff[1982] = 64'hffffa45affffa6a5;
    assign coff[1983] = 64'hffff8003fffffe61;
    assign coff[1984] = 64'hffff800afffffce8;
    assign coff[1985] = 64'hffffa355ffffa7b4;
    assign coff[1986] = 64'hffff8af6ffffcc2d;
    assign coff[1987] = 64'hffff8898ffffd1e3;
    assign coff[1988] = 64'hffff8319ffffe401;
    assign coff[1989] = 64'hffff93e3ffffbb7b;
    assign coff[1990] = 64'hffff9752ffffb656;
    assign coff[1991] = 64'hffff81e5ffffea12;
    assign coff[1992] = 64'hffff80f5fffff061;
    assign coff[1993] = 64'hffff9b1fffffb136;
    assign coff[1994] = 64'hffff909bffffc0f4;
    assign coff[1995] = 64'hffff84a6ffffddd0;
    assign coff[1996] = 64'hffff8672ffffd7e5;
    assign coff[1997] = 64'hffff8db0ffffc668;
    assign coff[1998] = 64'hffff9f0cffffac6e;
    assign coff[1999] = 64'hffff805afffff689;
    assign coff[2000] = 64'hffff8058fffff6a2;
    assign coff[2001] = 64'hffff9f1cffffac5b;
    assign coff[2002] = 64'hffff8da5ffffc67e;
    assign coff[2003] = 64'hffff867affffd7cd;
    assign coff[2004] = 64'hffff84a0ffffdde8;
    assign coff[2005] = 64'hffff90a7ffffc0de;
    assign coff[2006] = 64'hffff9b10ffffb14a;
    assign coff[2007] = 64'hffff80f8fffff048;
    assign coff[2008] = 64'hffff81e0ffffea2a;
    assign coff[2009] = 64'hffff9761ffffb642;
    assign coff[2010] = 64'hffff93d5ffffbb90;
    assign coff[2011] = 64'hffff831fffffe3e8;
    assign coff[2012] = 64'hffff888fffffd1fb;
    assign coff[2013] = 64'hffff8b00ffffcc16;
    assign coff[2014] = 64'hffffa343ffffa7c6;
    assign coff[2015] = 64'hffff800afffffccf;
    assign coff[2016] = 64'hffff8027fffff9c5;
    assign coff[2017] = 64'hffffa131ffffaa01;
    assign coff[2018] = 64'hffff8c45ffffc951;
    assign coff[2019] = 64'hffff8780ffffd4d5;
    assign coff[2020] = 64'hffff83d3ffffe0f2;
    assign coff[2021] = 64'hffff923cffffbe27;
    assign coff[2022] = 64'hffff9929ffffb3ca;
    assign coff[2023] = 64'hffff8165ffffed2c;
    assign coff[2024] = 64'hffff8161ffffed44;
    assign coff[2025] = 64'hffff9938ffffb3b6;
    assign coff[2026] = 64'hffff922fffffbe3d;
    assign coff[2027] = 64'hffff83d9ffffe0da;
    assign coff[2028] = 64'hffff8777ffffd4ed;
    assign coff[2029] = 64'hffff8c4fffffc93b;
    assign coff[2030] = 64'hffffa120ffffaa14;
    assign coff[2031] = 64'hffff8028fffff9ac;
    assign coff[2032] = 64'hffff809dfffff381;
    assign coff[2033] = 64'hffff9d16ffffaec2;
    assign coff[2034] = 64'hffff8f17ffffc3b4;
    assign coff[2035] = 64'hffff8587ffffdacc;
    assign coff[2036] = 64'hffff857fffffdae4;
    assign coff[2037] = 64'hffff8f23ffffc39e;
    assign coff[2038] = 64'hffff9d06ffffaed6;
    assign coff[2039] = 64'hffff809ffffff368;
    assign coff[2040] = 64'hffff8273ffffe714;
    assign coff[2041] = 64'hffff9599ffffb8d9;
    assign coff[2042] = 64'hffff958bffffb8ee;
    assign coff[2043] = 64'hffff8278ffffe6fb;
    assign coff[2044] = 64'hffff89baffffcf10;
    assign coff[2045] = 64'hffff89c3ffffcef9;
    assign coff[2046] = 64'hffffa575ffffa586;
    assign coff[2047] = 64'hffff8000fffffff3;




    always_ff @(posedge clk, negedge rst_n) begin
        if(~rst_n) begin
            data_o_col1 <= 'b0;
            data_o_col2 <= 'b0;
        end else begin
            if ((addr_col1 == 'd0 || addr_col1 == 'd1) && (valid == 1)) begin
                data_o_col1 <= coff[addr_col1];
                data_o_col2 <= 'b0;
            end else if(valid == 1) begin
                data_o_col1 <= coff[addr_col1];
                data_o_col2 <= coff[addr_col2];
            end begin
                data_o_col1 <= 'b0;
                data_o_col2 <= 'b0;
            end       
        end
    end


endmodule