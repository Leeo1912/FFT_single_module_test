// `timescale 1ns/1ps
module rom_3
(
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic                     valid,
    input  logic [10:0]              addr_i,
    output logic [255:0]              data_o
);

    logic [255:0] coff[2047:0];

    assign coff[0   ] = 256'h00007fff000000000000000000007fffffff80010000000000000000ffff8001;
    assign coff[1   ] = 256'hffffa57effffa57e00005a82ffffa57e00005a8200005a82ffffa57e00005a82;
    assign coff[2   ] = 256'h000030fcffff89be00007642000030fcffffcf0400007642ffff89beffffcf04;
    assign coff[3   ] = 256'hffff89be000030fcffffcf04ffff89be00007642ffffcf04000030fc00007642;
    assign coff[4   ] = 256'h00006a6effffb8e30000471d00006a6effff95920000471dffffb8e3ffff9592;
    assign coff[5   ] = 256'hffff8276ffffe707000018f9ffff827600007d8a000018f9ffffe70700007d8a;
    assign coff[6   ] = 256'hffffe707ffff827600007d8affffe707000018f900007d8affff8276000018f9;
    assign coff[7   ] = 256'hffffb8e300006a6effff9592ffffb8e30000471dffff959200006a6e0000471d;
    assign coff[8   ] = 256'h00007a7dffffdad80000252800007a7dffff858300002528ffffdad8ffff8583;
    assign coff[9   ] = 256'hffff8f1dffffc3a900003c57ffff8f1d000070e300003c57ffffc3a9000070e3;
    assign coff[10  ] = 256'h00000c8cffff809e00007f6200000c8cfffff37400007f62ffff809efffff374;
    assign coff[11  ] = 256'hffff9d0e00005134ffffaeccffff9d0e000062f2ffffaecc00005134000062f2;
    assign coff[12  ] = 256'h00005134ffff9d0e000062f200005134ffffaecc000062f2ffff9d0effffaecc;
    assign coff[13  ] = 256'hffff809e00000c8cfffff374ffff809e00007f62fffff37400000c8c00007f62;
    assign coff[14  ] = 256'hffffc3a9ffff8f1d000070e3ffffc3a900003c57000070e3ffff8f1d00003c57;
    assign coff[15  ] = 256'hffffdad800007a7dffff8583ffffdad800002528ffff858300007a7d00002528;
    assign coff[16  ] = 256'h00007e9dffffed38000012c800007e9dffff8163000012c8ffffed38ffff8163;
    assign coff[17  ] = 256'hffff9930ffffb3c000004c40ffff9930000066d000004c40ffffb3c0000066d0;
    assign coff[18  ] = 256'h00001f1affff83d600007c2a00001f1affffe0e600007c2affff83d6ffffe0e6;
    assign coff[19  ] = 256'hffff9236000041ceffffbe32ffff923600006dcaffffbe32000041ce00006dca;
    assign coff[20  ] = 256'h00005ed7ffffaa0a000055f600005ed7ffffa129000055f6ffffaa0affffa129;
    assign coff[21  ] = 256'hffff8027fffff9b800000648ffff802700007fd900000648fffff9b800007fd9;
    assign coff[22  ] = 256'hffffd4e1ffff877b00007885ffffd4e100002b1f00007885ffff877b00002b1f;
    assign coff[23  ] = 256'hffffc946000073b6ffff8c4affffc946000036baffff8c4a000073b6000036ba;
    assign coff[24  ] = 256'h000073b6ffffc946000036ba000073b6ffff8c4a000036baffffc946ffff8c4a;
    assign coff[25  ] = 256'hffff877bffffd4e100002b1fffff877b0000788500002b1fffffd4e100007885;
    assign coff[26  ] = 256'hfffff9b8ffff802700007fd9fffff9b80000064800007fd9ffff802700000648;
    assign coff[27  ] = 256'hffffaa0a00005ed7ffffa129ffffaa0a000055f6ffffa12900005ed7000055f6;
    assign coff[28  ] = 256'h000041ceffff923600006dca000041ceffffbe3200006dcaffff9236ffffbe32;
    assign coff[29  ] = 256'hffff83d600001f1affffe0e6ffff83d600007c2affffe0e600001f1a00007c2a;
    assign coff[30  ] = 256'hffffb3c0ffff9930000066d0ffffb3c000004c40000066d0ffff993000004c40;
    assign coff[31  ] = 256'hffffed3800007e9dffff8163ffffed38000012c8ffff816300007e9d000012c8;
    assign coff[32  ] = 256'h00007fa7fffff6950000096b00007fa7ffff80590000096bfffff695ffff8059;
    assign coff[33  ] = 256'hffff9f14ffffac650000539bffff9f14000060ec0000539bffffac65000060ec;
    assign coff[34  ] = 256'h00002827ffff86760000798a00002827ffffd7d90000798affff8676ffffd7d9;
    assign coff[35  ] = 256'hffff8dab0000398dffffc673ffff8dab00007255ffffc6730000398d00007255;
    assign coff[36  ] = 256'h000064e9ffffb14000004ec0000064e9ffff9b1700004ec0ffffb140ffff9b17;
    assign coff[37  ] = 256'hffff80f6fffff05500000fabffff80f600007f0a00000fabfffff05500007f0a;
    assign coff[38  ] = 256'hffffdddcffff84a300007b5dffffdddc0000222400007b5dffff84a300002224;
    assign coff[39  ] = 256'hffffc0e900006f5fffff90a1ffffc0e900003f17ffff90a100006f5f00003f17;
    assign coff[40  ] = 256'h0000776cffffd1ef00002e110000776cffff889400002e11ffffd1efffff8894;
    assign coff[41  ] = 256'hffff8afbffffcc21000033dfffff8afb00007505000033dfffffcc2100007505;
    assign coff[42  ] = 256'h00000324ffff800a00007ff600000324fffffcdc00007ff6ffff800afffffcdc;
    assign coff[43  ] = 256'hffffa34c00005843ffffa7bdffffa34c00005cb4ffffa7bd0000584300005cb4;
    assign coff[44  ] = 256'h000049b4ffff9759000068a7000049b4ffffb64c000068a7ffff9759ffffb64c;
    assign coff[45  ] = 256'hffff81e2000015e2ffffea1effff81e200007e1effffea1e000015e200007e1e;
    assign coff[46  ] = 256'hffffbb85ffff93dc00006c24ffffbb850000447b00006c24ffff93dc0000447b;
    assign coff[47  ] = 256'hffffe3f400007ce4ffff831cffffe3f400001c0cffff831c00007ce400001c0c;
    assign coff[48  ] = 256'h00007ce4ffffe3f400001c0c00007ce4ffff831c00001c0cffffe3f4ffff831c;
    assign coff[49  ] = 256'hffff93dcffffbb850000447bffff93dc00006c240000447bffffbb8500006c24;
    assign coff[50  ] = 256'h000015e2ffff81e200007e1e000015e2ffffea1e00007e1effff81e2ffffea1e;
    assign coff[51  ] = 256'hffff9759000049b4ffffb64cffff9759000068a7ffffb64c000049b4000068a7;
    assign coff[52  ] = 256'h00005843ffffa34c00005cb400005843ffffa7bd00005cb4ffffa34cffffa7bd;
    assign coff[53  ] = 256'hffff800a00000324fffffcdcffff800a00007ff6fffffcdc0000032400007ff6;
    assign coff[54  ] = 256'hffffcc21ffff8afb00007505ffffcc21000033df00007505ffff8afb000033df;
    assign coff[55  ] = 256'hffffd1ef0000776cffff8894ffffd1ef00002e11ffff88940000776c00002e11;
    assign coff[56  ] = 256'h00006f5fffffc0e900003f1700006f5fffff90a100003f17ffffc0e9ffff90a1;
    assign coff[57  ] = 256'hffff84a3ffffdddc00002224ffff84a300007b5d00002224ffffdddc00007b5d;
    assign coff[58  ] = 256'hfffff055ffff80f600007f0afffff05500000fab00007f0affff80f600000fab;
    assign coff[59  ] = 256'hffffb140000064e9ffff9b17ffffb14000004ec0ffff9b17000064e900004ec0;
    assign coff[60  ] = 256'h0000398dffff8dab000072550000398dffffc67300007255ffff8dabffffc673;
    assign coff[61  ] = 256'hffff867600002827ffffd7d9ffff86760000798affffd7d9000028270000798a;
    assign coff[62  ] = 256'hffffac65ffff9f14000060ecffffac650000539b000060ecffff9f140000539b;
    assign coff[63  ] = 256'hfffff69500007fa7ffff8059fffff6950000096bffff805900007fa70000096b;
    assign coff[64  ] = 256'h00007feafffffb4a000004b600007feaffff8016000004b6fffffb4affff8016;
    assign coff[65  ] = 256'hffffa238ffffa8e20000571effffa23800005dc80000571effffa8e200005dc8;
    assign coff[66  ] = 256'h00002c99ffff8805000077fb00002c99ffffd367000077fbffff8805ffffd367;
    assign coff[67  ] = 256'hffff8ba00000354effffcab2ffff8ba000007460ffffcab20000354e00007460;
    assign coff[68  ] = 256'h000067bdffffb50500004afb000067bdffff984300004afbffffb505ffff9843;
    assign coff[69  ] = 256'hffff81a0ffffebab00001455ffff81a000007e6000001455ffffebab00007e60;
    assign coff[70  ] = 256'hffffe26dffff837700007c89ffffe26d00001d9300007c89ffff837700001d93;
    assign coff[71  ] = 256'hffffbcda00006cf9ffff9307ffffbcda00004326ffff930700006cf900004326;
    assign coff[72  ] = 256'h0000790affffd65c000029a40000790affff86f6000029a4ffffd65cffff86f6;
    assign coff[73  ] = 256'hffff8cf8ffffc7db00003825ffff8cf80000730800003825ffffc7db00007308;
    assign coff[74  ] = 256'h000007d9ffff803e00007fc2000007d9fffff82700007fc2ffff803efffff827;
    assign coff[75  ] = 256'hffffa01c000054caffffab36ffffa01c00005fe4ffffab36000054ca00005fe4;
    assign coff[76  ] = 256'h00004d81ffff9a22000065de00004d81ffffb27f000065deffff9a22ffffb27f;
    assign coff[77  ] = 256'hffff812a0000113affffeec6ffff812a00007ed6ffffeec60000113a00007ed6;
    assign coff[78  ] = 256'hffffbf8cffff916900006e97ffffbf8c0000407400006e97ffff916900004074;
    assign coff[79  ] = 256'hffffdf6100007bc6ffff843affffdf610000209fffff843a00007bc60000209f;
    assign coff[80  ] = 256'h00007dd6ffffe8920000176e00007dd6ffff822a0000176effffe892ffff822a;
    assign coff[81  ] = 256'hffff9674ffffb7960000486affff96740000698c0000486affffb7960000698c;
    assign coff[82  ] = 256'h00001a83ffff82c600007d3a00001a83ffffe57d00007d3affff82c6ffffe57d;
    assign coff[83  ] = 256'hffff94b5000045cdffffba33ffff94b500006b4bffffba33000045cd00006b4b;
    assign coff[84  ] = 256'h00005b9dffffa69c0000596400005b9dffffa46300005964ffffa69cffffa463;
    assign coff[85  ] = 256'hffff8002fffffe6e00000192ffff800200007ffe00000192fffffe6e00007ffe;
    assign coff[86  ] = 256'hffffd079ffff8927000076d9ffffd07900002f87000076d9ffff892700002f87;
    assign coff[87  ] = 256'hffffcd92000075a6ffff8a5affffcd920000326effff8a5a000075a60000326e;
    assign coff[88  ] = 256'h0000719effffc50d00003af30000719effff8e6200003af3ffffc50dffff8e62;
    assign coff[89  ] = 256'hffff85faffffd958000026a8ffff85fa00007a06000026a8ffffd95800007a06;
    assign coff[90  ] = 256'hfffff505ffff807900007f87fffff50500000afb00007f87ffff807900000afb;
    assign coff[91  ] = 256'hffffad97000061f1ffff9e0fffffad9700005269ffff9e0f000061f100005269;
    assign coff[92  ] = 256'h00003db8ffff8fdd0000702300003db8ffffc24800007023ffff8fddffffc248;
    assign coff[93  ] = 256'hffff8511000023a7ffffdc59ffff851100007aefffffdc59000023a700007aef;
    assign coff[94  ] = 256'hffffb005ffff9c11000063efffffb00500004ffb000063efffff9c1100004ffb;
    assign coff[95  ] = 256'hfffff1e400007f38ffff80c8fffff1e400000e1cffff80c800007f3800000e1c;
    assign coff[96  ] = 256'h00007f38fffff1e400000e1c00007f38ffff80c800000e1cfffff1e4ffff80c8;
    assign coff[97  ] = 256'hffff9c11ffffb00500004ffbffff9c11000063ef00004ffbffffb005000063ef;
    assign coff[98  ] = 256'h000023a7ffff851100007aef000023a7ffffdc5900007aefffff8511ffffdc59;
    assign coff[99  ] = 256'hffff8fdd00003db8ffffc248ffff8fdd00007023ffffc24800003db800007023;
    assign coff[100 ] = 256'h000061f1ffffad9700005269000061f1ffff9e0f00005269ffffad97ffff9e0f;
    assign coff[101 ] = 256'hffff8079fffff50500000afbffff807900007f8700000afbfffff50500007f87;
    assign coff[102 ] = 256'hffffd958ffff85fa00007a06ffffd958000026a800007a06ffff85fa000026a8;
    assign coff[103 ] = 256'hffffc50d0000719effff8e62ffffc50d00003af3ffff8e620000719e00003af3;
    assign coff[104 ] = 256'h000075a6ffffcd920000326e000075a6ffff8a5a0000326effffcd92ffff8a5a;
    assign coff[105 ] = 256'hffff8927ffffd07900002f87ffff8927000076d900002f87ffffd079000076d9;
    assign coff[106 ] = 256'hfffffe6effff800200007ffefffffe6e0000019200007ffeffff800200000192;
    assign coff[107 ] = 256'hffffa69c00005b9dffffa463ffffa69c00005964ffffa46300005b9d00005964;
    assign coff[108 ] = 256'h000045cdffff94b500006b4b000045cdffffba3300006b4bffff94b5ffffba33;
    assign coff[109 ] = 256'hffff82c600001a83ffffe57dffff82c600007d3affffe57d00001a8300007d3a;
    assign coff[110 ] = 256'hffffb796ffff96740000698cffffb7960000486a0000698cffff96740000486a;
    assign coff[111 ] = 256'hffffe89200007dd6ffff822affffe8920000176effff822a00007dd60000176e;
    assign coff[112 ] = 256'h00007bc6ffffdf610000209f00007bc6ffff843a0000209fffffdf61ffff843a;
    assign coff[113 ] = 256'hffff9169ffffbf8c00004074ffff916900006e9700004074ffffbf8c00006e97;
    assign coff[114 ] = 256'h0000113affff812a00007ed60000113affffeec600007ed6ffff812affffeec6;
    assign coff[115 ] = 256'hffff9a2200004d81ffffb27fffff9a22000065deffffb27f00004d81000065de;
    assign coff[116 ] = 256'h000054caffffa01c00005fe4000054caffffab3600005fe4ffffa01cffffab36;
    assign coff[117 ] = 256'hffff803e000007d9fffff827ffff803e00007fc2fffff827000007d900007fc2;
    assign coff[118 ] = 256'hffffc7dbffff8cf800007308ffffc7db0000382500007308ffff8cf800003825;
    assign coff[119 ] = 256'hffffd65c0000790affff86f6ffffd65c000029a4ffff86f60000790a000029a4;
    assign coff[120 ] = 256'h00006cf9ffffbcda0000432600006cf9ffff930700004326ffffbcdaffff9307;
    assign coff[121 ] = 256'hffff8377ffffe26d00001d93ffff837700007c8900001d93ffffe26d00007c89;
    assign coff[122 ] = 256'hffffebabffff81a000007e60ffffebab0000145500007e60ffff81a000001455;
    assign coff[123 ] = 256'hffffb505000067bdffff9843ffffb50500004afbffff9843000067bd00004afb;
    assign coff[124 ] = 256'h0000354effff8ba0000074600000354effffcab200007460ffff8ba0ffffcab2;
    assign coff[125 ] = 256'hffff880500002c99ffffd367ffff8805000077fbffffd36700002c99000077fb;
    assign coff[126 ] = 256'hffffa8e2ffffa23800005dc8ffffa8e20000571e00005dc8ffffa2380000571e;
    assign coff[127 ] = 256'hfffffb4a00007feaffff8016fffffb4a000004b6ffff801600007fea000004b6;
    assign coff[128 ] = 256'h00007ffafffffda50000025b00007ffaffff80060000025bfffffda5ffff8006;
    assign coff[129 ] = 256'hffffa3d7ffffa72c000058d4ffffa3d700005c29000058d4ffffa72c00005c29;
    assign coff[130 ] = 256'h00002eccffff88dd0000772300002eccffffd13400007723ffff88ddffffd134;
    assign coff[131 ] = 256'hffff8aaa00003327ffffccd9ffff8aaa00007556ffffccd90000332700007556;
    assign coff[132 ] = 256'h0000691affffb6f10000490f0000691affff96e60000490fffffb6f1ffff96e6;
    assign coff[133 ] = 256'hffff8205ffffe958000016a8ffff820500007dfb000016a8ffffe95800007dfb;
    assign coff[134 ] = 256'hffffe4b9ffff82f100007d0fffffe4b900001b4700007d0fffff82f100001b47;
    assign coff[135 ] = 256'hffffbadc00006bb8ffff9448ffffbadc00004524ffff944800006bb800004524;
    assign coff[136 ] = 256'h000079c9ffffd89800002768000079c9ffff863700002768ffffd898ffff8637;
    assign coff[137 ] = 256'hffff8e06ffffc5c000003a40ffff8e06000071fa00003a40ffffc5c0000071fa;
    assign coff[138 ] = 256'h00000a33ffff806800007f9800000a33fffff5cd00007f98ffff8068fffff5cd;
    assign coff[139 ] = 256'hffff9e9100005303ffffacfdffff9e910000616fffffacfd000053030000616f;
    assign coff[140 ] = 256'h00004f5effff9b940000646c00004f5effffb0a20000646cffff9b94ffffb0a2;
    assign coff[141 ] = 256'hffff80de00000ee4fffff11cffff80de00007f22fffff11c00000ee400007f22;
    assign coff[142 ] = 256'hffffc198ffff903e00006fc2ffffc19800003e6800006fc2ffff903e00003e68;
    assign coff[143 ] = 256'hffffdd1b00007b27ffff84d9ffffdd1b000022e5ffff84d900007b27000022e5;
    assign coff[144 ] = 256'h00007e3fffffeae40000151c00007e3fffff81c10000151cffffeae4ffff81c1;
    assign coff[145 ] = 256'hffff97ceffffb5a800004a58ffff97ce0000683200004a58ffffb5a800006832;
    assign coff[146 ] = 256'h00001cd0ffff834900007cb700001cd0ffffe33000007cb7ffff8349ffffe330;
    assign coff[147 ] = 256'hffff9371000043d1ffffbc2fffff937100006c8fffffbc2f000043d100006c8f;
    assign coff[148 ] = 256'h00005d3effffa84f000057b100005d3effffa2c2000057b1ffffa84fffffa2c2;
    assign coff[149 ] = 256'hffff800ffffffc13000003edffff800f00007ff1000003edfffffc1300007ff1;
    assign coff[150 ] = 256'hffffd2abffff884c000077b4ffffd2ab00002d55000077b4ffff884c00002d55;
    assign coff[151 ] = 256'hffffcb69000074b3ffff8b4dffffcb6900003497ffff8b4d000074b300003497;
    assign coff[152 ] = 256'h000072afffffc727000038d9000072afffff8d51000038d9ffffc727ffff8d51;
    assign coff[153 ] = 256'hffff86b6ffffd71b000028e5ffff86b60000794a000028e5ffffd71b0000794a;
    assign coff[154 ] = 256'hfffff75effff804b00007fb5fffff75e000008a200007fb5ffff804b000008a2;
    assign coff[155 ] = 256'hffffabcd00006068ffff9f98ffffabcd00005433ffff9f980000606800005433;
    assign coff[156 ] = 256'h00003fc6ffff910500006efb00003fc6ffffc03a00006efbffff9105ffffc03a;
    assign coff[157 ] = 256'hffff846e00002162ffffde9effff846e00007b92ffffde9e0000216200007b92;
    assign coff[158 ] = 256'hffffb1dfffff9a9c00006564ffffb1df00004e2100006564ffff9a9c00004e21;
    assign coff[159 ] = 256'hffffef8d00007ef0ffff8110ffffef8d00001073ffff811000007ef000001073;
    assign coff[160 ] = 256'h00007f75fffff43c00000bc400007f75ffff808b00000bc4fffff43cffff808b;
    assign coff[161 ] = 256'hffff9d8effffae31000051cfffff9d8e00006272000051cfffffae3100006272;
    assign coff[162 ] = 256'h000025e8ffff85be00007a42000025e8ffffda1800007a42ffff85beffffda18;
    assign coff[163 ] = 256'hffff8ebf00003ba5ffffc45bffff8ebf00007141ffffc45b00003ba500007141;
    assign coff[164 ] = 256'h00006371ffffaf680000509800006371ffff9c8f00005098ffffaf68ffff9c8f;
    assign coff[165 ] = 256'hffff80b2fffff2ac00000d54ffff80b200007f4e00000d54fffff2ac00007f4e;
    assign coff[166 ] = 256'hffffdb99ffff854900007ab7ffffdb990000246700007ab7ffff854900002467;
    assign coff[167 ] = 256'hffffc2f800007083ffff8f7dffffc2f800003d08ffff8f7d0000708300003d08;
    assign coff[168 ] = 256'h0000768effffcfbe000030420000768effff897200003042ffffcfbeffff8972;
    assign coff[169 ] = 256'hffff8a0cffffce4b000031b5ffff8a0c000075f4000031b5ffffce4b000075f4;
    assign coff[170 ] = 256'h000000c9ffff800100007fff000000c9ffffff3700007fffffff8001ffffff37;
    assign coff[171 ] = 256'hffffa4f0000059f4ffffa60cffffa4f000005b10ffffa60c000059f400005b10;
    assign coff[172 ] = 256'h000047c4ffff9603000069fd000047c4ffffb83c000069fdffff9603ffffb83c;
    assign coff[173 ] = 256'hffff824f00001833ffffe7cdffff824f00007db1ffffe7cd0000183300007db1;
    assign coff[174 ] = 256'hffffb98bffff952300006addffffb98b0000467500006addffff952300004675;
    assign coff[175 ] = 256'hffffe64200007d63ffff829dffffe642000019beffff829d00007d63000019be;
    assign coff[176 ] = 256'h00007c5affffe1a900001e5700007c5affff83a600001e57ffffe1a9ffff83a6;
    assign coff[177 ] = 256'hffff929effffbd860000427affff929e00006d620000427affffbd8600006d62;
    assign coff[178 ] = 256'h0000138fffff818100007e7f0000138fffffec7100007e7fffff8181ffffec71;
    assign coff[179 ] = 256'hffff98b900004b9effffb462ffff98b900006747ffffb46200004b9e00006747;
    assign coff[180 ] = 256'h0000568affffa1b000005e500000568affffa97600005e50ffffa1b0ffffa976;
    assign coff[181 ] = 256'hffff801e0000057ffffffa81ffff801e00007fe2fffffa810000057f00007fe2;
    assign coff[182 ] = 256'hffffc9fcffff8bf50000740bffffc9fc000036040000740bffff8bf500003604;
    assign coff[183 ] = 256'hffffd42400007840ffff87c0ffffd42400002bdcffff87c00000784000002bdc;
    assign coff[184 ] = 256'h00006e31ffffbedf0000412100006e31ffff91cf00004121ffffbedfffff91cf;
    assign coff[185 ] = 256'hffff8407ffffe02300001fddffff840700007bf900001fddffffe02300007bf9;
    assign coff[186 ] = 256'hffffedffffff814600007ebaffffedff0000120100007ebaffff814600001201;
    assign coff[187 ] = 256'hffffb31f00006657ffff99a9ffffb31f00004ce1ffff99a90000665700004ce1;
    assign coff[188 ] = 256'h00003770ffff8ca10000735f00003770ffffc8900000735fffff8ca1ffffc890;
    assign coff[189 ] = 256'hffff873800002a62ffffd59effff8738000078c8ffffd59e00002a62000078c8;
    assign coff[190 ] = 256'hffffaaa0ffffa0a200005f5effffaaa00000556000005f5effffa0a200005560;
    assign coff[191 ] = 256'hfffff8ef00007fceffff8032fffff8ef00000711ffff803200007fce00000711;
    assign coff[192 ] = 256'h00007fcefffff8ef0000071100007fceffff803200000711fffff8efffff8032;
    assign coff[193 ] = 256'hffffa0a2ffffaaa000005560ffffa0a200005f5e00005560ffffaaa000005f5e;
    assign coff[194 ] = 256'h00002a62ffff8738000078c800002a62ffffd59e000078c8ffff8738ffffd59e;
    assign coff[195 ] = 256'hffff8ca100003770ffffc890ffff8ca10000735fffffc890000037700000735f;
    assign coff[196 ] = 256'h00006657ffffb31f00004ce100006657ffff99a900004ce1ffffb31fffff99a9;
    assign coff[197 ] = 256'hffff8146ffffedff00001201ffff814600007eba00001201ffffedff00007eba;
    assign coff[198 ] = 256'hffffe023ffff840700007bf9ffffe02300001fdd00007bf9ffff840700001fdd;
    assign coff[199 ] = 256'hffffbedf00006e31ffff91cfffffbedf00004121ffff91cf00006e3100004121;
    assign coff[200 ] = 256'h00007840ffffd42400002bdc00007840ffff87c000002bdcffffd424ffff87c0;
    assign coff[201 ] = 256'hffff8bf5ffffc9fc00003604ffff8bf50000740b00003604ffffc9fc0000740b;
    assign coff[202 ] = 256'h0000057fffff801e00007fe20000057ffffffa8100007fe2ffff801efffffa81;
    assign coff[203 ] = 256'hffffa1b00000568affffa976ffffa1b000005e50ffffa9760000568a00005e50;
    assign coff[204 ] = 256'h00004b9effff98b90000674700004b9effffb46200006747ffff98b9ffffb462;
    assign coff[205 ] = 256'hffff81810000138fffffec71ffff818100007e7fffffec710000138f00007e7f;
    assign coff[206 ] = 256'hffffbd86ffff929e00006d62ffffbd860000427a00006d62ffff929e0000427a;
    assign coff[207 ] = 256'hffffe1a900007c5affff83a6ffffe1a900001e57ffff83a600007c5a00001e57;
    assign coff[208 ] = 256'h00007d63ffffe642000019be00007d63ffff829d000019beffffe642ffff829d;
    assign coff[209 ] = 256'hffff9523ffffb98b00004675ffff952300006add00004675ffffb98b00006add;
    assign coff[210 ] = 256'h00001833ffff824f00007db100001833ffffe7cd00007db1ffff824fffffe7cd;
    assign coff[211 ] = 256'hffff9603000047c4ffffb83cffff9603000069fdffffb83c000047c4000069fd;
    assign coff[212 ] = 256'h000059f4ffffa4f000005b10000059f4ffffa60c00005b10ffffa4f0ffffa60c;
    assign coff[213 ] = 256'hffff8001000000c9ffffff37ffff800100007fffffffff37000000c900007fff;
    assign coff[214 ] = 256'hffffce4bffff8a0c000075f4ffffce4b000031b5000075f4ffff8a0c000031b5;
    assign coff[215 ] = 256'hffffcfbe0000768effff8972ffffcfbe00003042ffff89720000768e00003042;
    assign coff[216 ] = 256'h00007083ffffc2f800003d0800007083ffff8f7d00003d08ffffc2f8ffff8f7d;
    assign coff[217 ] = 256'hffff8549ffffdb9900002467ffff854900007ab700002467ffffdb9900007ab7;
    assign coff[218 ] = 256'hfffff2acffff80b200007f4efffff2ac00000d5400007f4effff80b200000d54;
    assign coff[219 ] = 256'hffffaf6800006371ffff9c8fffffaf6800005098ffff9c8f0000637100005098;
    assign coff[220 ] = 256'h00003ba5ffff8ebf0000714100003ba5ffffc45b00007141ffff8ebfffffc45b;
    assign coff[221 ] = 256'hffff85be000025e8ffffda18ffff85be00007a42ffffda18000025e800007a42;
    assign coff[222 ] = 256'hffffae31ffff9d8e00006272ffffae31000051cf00006272ffff9d8e000051cf;
    assign coff[223 ] = 256'hfffff43c00007f75ffff808bfffff43c00000bc4ffff808b00007f7500000bc4;
    assign coff[224 ] = 256'h00007ef0ffffef8d0000107300007ef0ffff811000001073ffffef8dffff8110;
    assign coff[225 ] = 256'hffff9a9cffffb1df00004e21ffff9a9c0000656400004e21ffffb1df00006564;
    assign coff[226 ] = 256'h00002162ffff846e00007b9200002162ffffde9e00007b92ffff846effffde9e;
    assign coff[227 ] = 256'hffff910500003fc6ffffc03affff910500006efbffffc03a00003fc600006efb;
    assign coff[228 ] = 256'h00006068ffffabcd0000543300006068ffff9f9800005433ffffabcdffff9f98;
    assign coff[229 ] = 256'hffff804bfffff75e000008a2ffff804b00007fb5000008a2fffff75e00007fb5;
    assign coff[230 ] = 256'hffffd71bffff86b60000794affffd71b000028e50000794affff86b6000028e5;
    assign coff[231 ] = 256'hffffc727000072afffff8d51ffffc727000038d9ffff8d51000072af000038d9;
    assign coff[232 ] = 256'h000074b3ffffcb6900003497000074b3ffff8b4d00003497ffffcb69ffff8b4d;
    assign coff[233 ] = 256'hffff884cffffd2ab00002d55ffff884c000077b400002d55ffffd2ab000077b4;
    assign coff[234 ] = 256'hfffffc13ffff800f00007ff1fffffc13000003ed00007ff1ffff800f000003ed;
    assign coff[235 ] = 256'hffffa84f00005d3effffa2c2ffffa84f000057b1ffffa2c200005d3e000057b1;
    assign coff[236 ] = 256'h000043d1ffff937100006c8f000043d1ffffbc2f00006c8fffff9371ffffbc2f;
    assign coff[237 ] = 256'hffff834900001cd0ffffe330ffff834900007cb7ffffe33000001cd000007cb7;
    assign coff[238 ] = 256'hffffb5a8ffff97ce00006832ffffb5a800004a5800006832ffff97ce00004a58;
    assign coff[239 ] = 256'hffffeae400007e3fffff81c1ffffeae40000151cffff81c100007e3f0000151c;
    assign coff[240 ] = 256'h00007b27ffffdd1b000022e500007b27ffff84d9000022e5ffffdd1bffff84d9;
    assign coff[241 ] = 256'hffff903effffc19800003e68ffff903e00006fc200003e68ffffc19800006fc2;
    assign coff[242 ] = 256'h00000ee4ffff80de00007f2200000ee4fffff11c00007f22ffff80defffff11c;
    assign coff[243 ] = 256'hffff9b9400004f5effffb0a2ffff9b940000646cffffb0a200004f5e0000646c;
    assign coff[244 ] = 256'h00005303ffff9e910000616f00005303ffffacfd0000616fffff9e91ffffacfd;
    assign coff[245 ] = 256'hffff806800000a33fffff5cdffff806800007f98fffff5cd00000a3300007f98;
    assign coff[246 ] = 256'hffffc5c0ffff8e06000071faffffc5c000003a40000071faffff8e0600003a40;
    assign coff[247 ] = 256'hffffd898000079c9ffff8637ffffd89800002768ffff8637000079c900002768;
    assign coff[248 ] = 256'h00006bb8ffffbadc0000452400006bb8ffff944800004524ffffbadcffff9448;
    assign coff[249 ] = 256'hffff82f1ffffe4b900001b47ffff82f100007d0f00001b47ffffe4b900007d0f;
    assign coff[250 ] = 256'hffffe958ffff820500007dfbffffe958000016a800007dfbffff8205000016a8;
    assign coff[251 ] = 256'hffffb6f10000691affff96e6ffffb6f10000490fffff96e60000691a0000490f;
    assign coff[252 ] = 256'h00003327ffff8aaa0000755600003327ffffccd900007556ffff8aaaffffccd9;
    assign coff[253 ] = 256'hffff88dd00002eccffffd134ffff88dd00007723ffffd13400002ecc00007723;
    assign coff[254 ] = 256'hffffa72cffffa3d700005c29ffffa72c000058d400005c29ffffa3d7000058d4;
    assign coff[255 ] = 256'hfffffda500007ffaffff8006fffffda50000025bffff800600007ffa0000025b;
    assign coff[256 ] = 256'h00007ffffffffed20000012e00007fffffff80010000012efffffed2ffff8001;
    assign coff[257 ] = 256'hffffa4a9ffffa654000059acffffa4a900005b57000059acffffa65400005b57;
    assign coff[258 ] = 256'h00002fe5ffff894c000076b400002fe5ffffd01b000076b4ffff894cffffd01b;
    assign coff[259 ] = 256'hffff8a3300003212ffffcdeeffff8a33000075cdffffcdee00003212000075cd;
    assign coff[260 ] = 256'h000069c5ffffb7e900004817000069c5ffff963b00004817ffffb7e9ffff963b;
    assign coff[261 ] = 256'hffff823cffffe82f000017d1ffff823c00007dc4000017d1ffffe82f00007dc4;
    assign coff[262 ] = 256'hffffe5e0ffff82b200007d4effffe5e000001a2000007d4effff82b200001a20;
    assign coff[263 ] = 256'hffffb9df00006b14ffff94ecffffb9df00004621ffff94ec00006b1400004621;
    assign coff[264 ] = 256'h00007a24ffffd9b80000264800007a24ffff85dc00002648ffffd9b8ffff85dc;
    assign coff[265 ] = 256'hffff8e90ffffc4b400003b4cffff8e900000717000003b4cffffc4b400007170;
    assign coff[266 ] = 256'h00000b60ffff808200007f7e00000b60fffff4a000007f7effff8082fffff4a0;
    assign coff[267 ] = 256'hffff9dce0000521cffffade4ffff9dce00006232ffffade40000521c00006232;
    assign coff[268 ] = 256'h0000504affff9c50000063b00000504affffafb6000063b0ffff9c50ffffafb6;
    assign coff[269 ] = 256'hffff80bd00000db8fffff248ffff80bd00007f43fffff24800000db800007f43;
    assign coff[270 ] = 256'hffffc2a0ffff8fad00007053ffffc2a000003d6000007053ffff8fad00003d60;
    assign coff[271 ] = 256'hffffdbf900007ad3ffff852dffffdbf900002407ffff852d00007ad300002407;
    assign coff[272 ] = 256'h00007e70ffffec0e000013f200007e70ffff8190000013f2ffffec0effff8190;
    assign coff[273 ] = 256'hffff987effffb4b300004b4dffff987e0000678200004b4dffffb4b300006782;
    assign coff[274 ] = 256'h00001df5ffff838e00007c7200001df5ffffe20b00007c72ffff838effffe20b;
    assign coff[275 ] = 256'hffff92d2000042d0ffffbd30ffff92d200006d2effffbd30000042d000006d2e;
    assign coff[276 ] = 256'h00005e0cffffa92c000056d400005e0cffffa1f4000056d4ffffa92cffffa1f4;
    assign coff[277 ] = 256'hffff801afffffae50000051bffff801a00007fe60000051bfffffae500007fe6;
    assign coff[278 ] = 256'hffffd3c5ffff87e20000781effffd3c500002c3b0000781effff87e200002c3b;
    assign coff[279 ] = 256'hffffca5700007436ffff8bcaffffca57000035a9ffff8bca00007436000035a9;
    assign coff[280 ] = 256'h00007334ffffc836000037ca00007334ffff8ccc000037caffffc836ffff8ccc;
    assign coff[281 ] = 256'hffff8717ffffd5fd00002a03ffff8717000078e900002a03ffffd5fd000078e9;
    assign coff[282 ] = 256'hfffff88bffff803800007fc8fffff88b0000077500007fc8ffff803800000775;
    assign coff[283 ] = 256'hffffaaeb00005fa1ffffa05fffffaaeb00005515ffffa05f00005fa100005515;
    assign coff[284 ] = 256'h000040cbffff919c00006e64000040cbffffbf3500006e64ffff919cffffbf35;
    assign coff[285 ] = 256'hffff84210000203effffdfc2ffff842100007bdfffffdfc20000203e00007bdf;
    assign coff[286 ] = 256'hffffb2cfffff99e50000661bffffb2cf00004d310000661bffff99e500004d31;
    assign coff[287 ] = 256'hffffee6200007ec8ffff8138ffffee620000119effff813800007ec80000119e;
    assign coff[288 ] = 256'h00007f90fffff56900000a9700007f90ffff807000000a97fffff569ffff8070;
    assign coff[289 ] = 256'hffff9e50ffffad4a000052b6ffff9e50000061b0000052b6ffffad4a000061b0;
    assign coff[290 ] = 256'h00002708ffff8619000079e700002708ffffd8f8000079e7ffff8619ffffd8f8;
    assign coff[291 ] = 256'hffff8e3400003a9affffc566ffff8e34000071ccffffc56600003a9a000071cc;
    assign coff[292 ] = 256'h0000642effffb05300004fad0000642effff9bd200004fadffffb053ffff9bd2;
    assign coff[293 ] = 256'hffff80d3fffff18000000e80ffff80d300007f2d00000e80fffff18000007f2d;
    assign coff[294 ] = 256'hffffdcbaffff84f500007b0bffffdcba0000234600007b0bffff84f500002346;
    assign coff[295 ] = 256'hffffc1f000006ff2ffff900effffc1f000003e10ffff900e00006ff200003e10;
    assign coff[296 ] = 256'h000076feffffd0d600002f2a000076feffff890200002f2affffd0d6ffff8902;
    assign coff[297 ] = 256'hffff8a82ffffcd35000032cbffff8a820000757e000032cbffffcd350000757e;
    assign coff[298 ] = 256'h000001f7ffff800400007ffc000001f7fffffe0900007ffcffff8004fffffe09;
    assign coff[299 ] = 256'hffffa41d0000591cffffa6e4ffffa41d00005be3ffffa6e40000591c00005be3;
    assign coff[300 ] = 256'h000048bdffff96ad00006953000048bdffffb74300006953ffff96adffffb743;
    assign coff[301 ] = 256'hffff82170000170bffffe8f5ffff821700007de9ffffe8f50000170b00007de9;
    assign coff[302 ] = 256'hffffba87ffff947e00006b82ffffba870000457900006b82ffff947e00004579;
    assign coff[303 ] = 256'hffffe51b00007d25ffff82dbffffe51b00001ae5ffff82db00007d2500001ae5;
    assign coff[304 ] = 256'h00007ca0ffffe2cf00001d3100007ca0ffff836000001d31ffffe2cfffff8360;
    assign coff[305 ] = 256'hffff933cffffbc850000437bffff933c00006cc40000437bffffbc8500006cc4;
    assign coff[306 ] = 256'h000014b9ffff81b000007e50000014b9ffffeb4700007e50ffff81b0ffffeb47;
    assign coff[307 ] = 256'hffff980800004aaaffffb556ffff9808000067f8ffffb55600004aaa000067f8;
    assign coff[308 ] = 256'h00005767ffffa27d00005d8300005767ffffa89900005d83ffffa27dffffa899;
    assign coff[309 ] = 256'hffff801300000452fffffbaeffff801300007fedfffffbae0000045200007fed;
    assign coff[310 ] = 256'hffffcb0effff8b7700007489ffffcb0e000034f200007489ffff8b77000034f2;
    assign coff[311 ] = 256'hffffd309000077d8ffff8828ffffd30900002cf7ffff8828000077d800002cf7;
    assign coff[312 ] = 256'h00006ec9ffffbfe30000401d00006ec9ffff91370000401dffffbfe3ffff9137;
    assign coff[313 ] = 256'hffff8454ffffdeff00002101ffff845400007bac00002101ffffdeff00007bac;
    assign coff[314 ] = 256'hffffef2affff811d00007ee3ffffef2a000010d600007ee3ffff811d000010d6;
    assign coff[315 ] = 256'hffffb22f000065a1ffff9a5fffffb22f00004dd1ffff9a5f000065a100004dd1;
    assign coff[316 ] = 256'h0000387fffff8d24000072dc0000387fffffc781000072dcffff8d24ffffc781;
    assign coff[317 ] = 256'hffff86d600002945ffffd6bbffff86d60000792affffd6bb000029450000792a;
    assign coff[318 ] = 256'hffffab81ffff9fda00006026ffffab810000547f00006026ffff9fda0000547f;
    assign coff[319 ] = 256'hfffff7c200007fbcffff8044fffff7c20000083effff804400007fbc0000083e;
    assign coff[320 ] = 256'h00007fddfffffa1d000005e300007fddffff8023000005e3fffffa1dffff8023;
    assign coff[321 ] = 256'hffffa16cffffa9c000005640ffffa16c00005e9400005640ffffa9c000005e94;
    assign coff[322 ] = 256'h00002b7effff879d0000786300002b7effffd48200007863ffff879dffffd482;
    assign coff[323 ] = 256'hffff8c1f0000365fffffc9a1ffff8c1f000073e1ffffc9a10000365f000073e1;
    assign coff[324 ] = 256'h0000670bffffb41100004bef0000670bffff98f500004befffffb411ffff98f5;
    assign coff[325 ] = 256'hffff8172ffffecd50000132bffff817200007e8e0000132bffffecd500007e8e;
    assign coff[326 ] = 256'hffffe148ffff83be00007c42ffffe14800001eb800007c42ffff83be00001eb8;
    assign coff[327 ] = 256'hffffbddc00006d96ffff926affffbddc00004224ffff926a00006d9600004224;
    assign coff[328 ] = 256'h000078a6ffffd53f00002ac1000078a6ffff875a00002ac1ffffd53fffff875a;
    assign coff[329 ] = 256'hffff8c75ffffc8eb00003715ffff8c750000738b00003715ffffc8eb0000738b;
    assign coff[330 ] = 256'h000006acffff802d00007fd3000006acfffff95400007fd3ffff802dfffff954;
    assign coff[331 ] = 256'hffffa0e5000055abffffaa55ffffa0e500005f1bffffaa55000055ab00005f1b;
    assign coff[332 ] = 256'h00004c91ffff996d0000669300004c91ffffb36f00006693ffff996dffffb36f;
    assign coff[333 ] = 256'hffff815400001265ffffed9bffff815400007eacffffed9b0000126500007eac;
    assign coff[334 ] = 256'hffffbe88ffff920200006dfeffffbe880000417800006dfeffff920200004178;
    assign coff[335 ] = 256'hffffe08500007c11ffff83efffffe08500001f7bffff83ef00007c1100001f7b;
    assign coff[336 ] = 256'h00007d9effffe76a0000189600007d9effff826200001896ffffe76affff8262;
    assign coff[337 ] = 256'hffff95caffffb89000004770ffff95ca00006a3600004770ffffb89000006a36;
    assign coff[338 ] = 256'h0000195bffff828900007d770000195bffffe6a500007d77ffff8289ffffe6a5;
    assign coff[339 ] = 256'hffff955b000046c9ffffb937ffff955b00006aa5ffffb937000046c900006aa5;
    assign coff[340 ] = 256'h00005ac9ffffa5c500005a3b00005ac9ffffa53700005a3bffffa5c5ffffa537;
    assign coff[341 ] = 256'hffff8001ffffff9b00000065ffff800100007fff00000065ffffff9b00007fff;
    assign coff[342 ] = 256'hffffcf61ffff899800007668ffffcf610000309f00007668ffff89980000309f;
    assign coff[343 ] = 256'hffffcea70000761bffff89e5ffffcea700003159ffff89e50000761b00003159;
    assign coff[344 ] = 256'h00007112ffffc40200003bfe00007112ffff8eee00003bfeffffc402ffff8eee;
    assign coff[345 ] = 256'hffff85a0ffffda7800002588ffff85a000007a6000002588ffffda7800007a60;
    assign coff[346 ] = 256'hfffff3d8ffff809400007f6cfffff3d800000c2800007f6cffff809400000c28;
    assign coff[347 ] = 256'hffffae7f000062b2ffff9d4effffae7f00005181ffff9d4e000062b200005181;
    assign coff[348 ] = 256'h00003cafffff8f4d000070b300003cafffffc351000070b3ffff8f4dffffc351;
    assign coff[349 ] = 256'hffff8566000024c8ffffdb38ffff856600007a9affffdb38000024c800007a9a;
    assign coff[350 ] = 256'hffffaf1affff9cce00006332ffffaf1a000050e600006332ffff9cce000050e6;
    assign coff[351 ] = 256'hfffff31000007f58ffff80a8fffff31000000cf0ffff80a800007f5800000cf0;
    assign coff[352 ] = 256'h00007f16fffff0b900000f4700007f16ffff80ea00000f47fffff0b9ffff80ea;
    assign coff[353 ] = 256'hffff9b55ffffb0f100004f0fffff9b55000064ab00004f0fffffb0f1000064ab;
    assign coff[354 ] = 256'h00002284ffff84be00007b4200002284ffffdd7c00007b42ffff84beffffdd7c;
    assign coff[355 ] = 256'hffff907000003ec0ffffc140ffff907000006f90ffffc14000003ec000006f90;
    assign coff[356 ] = 256'h0000612effffacb10000534f0000612effff9ed20000534fffffacb1ffff9ed2;
    assign coff[357 ] = 256'hffff8060fffff631000009cfffff806000007fa0000009cffffff63100007fa0;
    assign coff[358 ] = 256'hffffd839ffff8656000079aaffffd839000027c7000079aaffff8656000027c7;
    assign coff[359 ] = 256'hffffc61900007228ffff8dd8ffffc619000039e7ffff8dd800007228000039e7;
    assign coff[360 ] = 256'h0000752dffffcc7d000033830000752dffff8ad300003383ffffcc7dffff8ad3;
    assign coff[361 ] = 256'hffff88b8ffffd19100002e6fffff88b80000774800002e6fffffd19100007748;
    assign coff[362 ] = 256'hfffffd40ffff800800007ff8fffffd40000002c000007ff8ffff8008000002c0;
    assign coff[363 ] = 256'hffffa77400005c6fffffa391ffffa7740000588cffffa39100005c6f0000588c;
    assign coff[364 ] = 256'h000044d0ffff941200006bee000044d0ffffbb3000006beeffff9412ffffbb30;
    assign coff[365 ] = 256'hffff830600001ba9ffffe457ffff830600007cfaffffe45700001ba900007cfa;
    assign coff[366 ] = 256'hffffb69effff9720000068e0ffffb69e00004962000068e0ffff972000004962;
    assign coff[367 ] = 256'hffffe9bb00007e0cffff81f4ffffe9bb00001645ffff81f400007e0c00001645;
    assign coff[368 ] = 256'h00007b78ffffde3d000021c300007b78ffff8488000021c3ffffde3dffff8488;
    assign coff[369 ] = 256'hffff90d3ffffc09100003f6fffff90d300006f2d00003f6fffffc09100006f2d;
    assign coff[370 ] = 256'h0000100fffff810300007efd0000100fffffeff100007efdffff8103ffffeff1;
    assign coff[371 ] = 256'hffff9ada00004e71ffffb18fffff9ada00006526ffffb18f00004e7100006526;
    assign coff[372 ] = 256'h000053e7ffff9f56000060aa000053e7ffffac19000060aaffff9f56ffffac19;
    assign coff[373 ] = 256'hffff805200000906fffff6faffff805200007faefffff6fa0000090600007fae;
    assign coff[374 ] = 256'hffffc6cdffff8d7e00007282ffffc6cd0000393300007282ffff8d7e00003933;
    assign coff[375 ] = 256'hffffd77a0000796affff8696ffffd77a00002886ffff86960000796a00002886;
    assign coff[376 ] = 256'h00006c5affffbbda0000442600006c5affff93a600004426ffffbbdaffff93a6;
    assign coff[377 ] = 256'hffff8332ffffe39200001c6effff833200007cce00001c6effffe39200007cce;
    assign coff[378 ] = 256'hffffea81ffff81d100007e2fffffea810000157f00007e2fffff81d10000157f;
    assign coff[379 ] = 256'hffffb5fa0000686dffff9793ffffb5fa00004a06ffff97930000686d00004a06;
    assign coff[380 ] = 256'h0000343bffff8b24000074dc0000343bffffcbc5000074dcffff8b24ffffcbc5;
    assign coff[381 ] = 256'hffff887000002db3ffffd24dffff887000007790ffffd24d00002db300007790;
    assign coff[382 ] = 256'hffffa806ffffa30700005cf9ffffa806000057fa00005cf9ffffa307000057fa;
    assign coff[383 ] = 256'hfffffc7700007ff4ffff800cfffffc7700000389ffff800c00007ff400000389;
    assign coff[384 ] = 256'h00007ff4fffffc770000038900007ff4ffff800c00000389fffffc77ffff800c;
    assign coff[385 ] = 256'hffffa307ffffa806000057faffffa30700005cf9000057faffffa80600005cf9;
    assign coff[386 ] = 256'h00002db3ffff88700000779000002db3ffffd24d00007790ffff8870ffffd24d;
    assign coff[387 ] = 256'hffff8b240000343bffffcbc5ffff8b24000074dcffffcbc50000343b000074dc;
    assign coff[388 ] = 256'h0000686dffffb5fa00004a060000686dffff979300004a06ffffb5faffff9793;
    assign coff[389 ] = 256'hffff81d1ffffea810000157fffff81d100007e2f0000157fffffea8100007e2f;
    assign coff[390 ] = 256'hffffe392ffff833200007cceffffe39200001c6e00007cceffff833200001c6e;
    assign coff[391 ] = 256'hffffbbda00006c5affff93a6ffffbbda00004426ffff93a600006c5a00004426;
    assign coff[392 ] = 256'h0000796affffd77a000028860000796affff869600002886ffffd77affff8696;
    assign coff[393 ] = 256'hffff8d7effffc6cd00003933ffff8d7e0000728200003933ffffc6cd00007282;
    assign coff[394 ] = 256'h00000906ffff805200007fae00000906fffff6fa00007faeffff8052fffff6fa;
    assign coff[395 ] = 256'hffff9f56000053e7ffffac19ffff9f56000060aaffffac19000053e7000060aa;
    assign coff[396 ] = 256'h00004e71ffff9ada0000652600004e71ffffb18f00006526ffff9adaffffb18f;
    assign coff[397 ] = 256'hffff81030000100fffffeff1ffff810300007efdffffeff10000100f00007efd;
    assign coff[398 ] = 256'hffffc091ffff90d300006f2dffffc09100003f6f00006f2dffff90d300003f6f;
    assign coff[399 ] = 256'hffffde3d00007b78ffff8488ffffde3d000021c3ffff848800007b78000021c3;
    assign coff[400 ] = 256'h00007e0cffffe9bb0000164500007e0cffff81f400001645ffffe9bbffff81f4;
    assign coff[401 ] = 256'hffff9720ffffb69e00004962ffff9720000068e000004962ffffb69e000068e0;
    assign coff[402 ] = 256'h00001ba9ffff830600007cfa00001ba9ffffe45700007cfaffff8306ffffe457;
    assign coff[403 ] = 256'hffff9412000044d0ffffbb30ffff941200006beeffffbb30000044d000006bee;
    assign coff[404 ] = 256'h00005c6fffffa7740000588c00005c6fffffa3910000588cffffa774ffffa391;
    assign coff[405 ] = 256'hffff8008fffffd40000002c0ffff800800007ff8000002c0fffffd4000007ff8;
    assign coff[406 ] = 256'hffffd191ffff88b800007748ffffd19100002e6f00007748ffff88b800002e6f;
    assign coff[407 ] = 256'hffffcc7d0000752dffff8ad3ffffcc7d00003383ffff8ad30000752d00003383;
    assign coff[408 ] = 256'h00007228ffffc619000039e700007228ffff8dd8000039e7ffffc619ffff8dd8;
    assign coff[409 ] = 256'hffff8656ffffd839000027c7ffff8656000079aa000027c7ffffd839000079aa;
    assign coff[410 ] = 256'hfffff631ffff806000007fa0fffff631000009cf00007fa0ffff8060000009cf;
    assign coff[411 ] = 256'hffffacb10000612effff9ed2ffffacb10000534fffff9ed20000612e0000534f;
    assign coff[412 ] = 256'h00003ec0ffff907000006f9000003ec0ffffc14000006f90ffff9070ffffc140;
    assign coff[413 ] = 256'hffff84be00002284ffffdd7cffff84be00007b42ffffdd7c0000228400007b42;
    assign coff[414 ] = 256'hffffb0f1ffff9b55000064abffffb0f100004f0f000064abffff9b5500004f0f;
    assign coff[415 ] = 256'hfffff0b900007f16ffff80eafffff0b900000f47ffff80ea00007f1600000f47;
    assign coff[416 ] = 256'h00007f58fffff31000000cf000007f58ffff80a800000cf0fffff310ffff80a8;
    assign coff[417 ] = 256'hffff9cceffffaf1a000050e6ffff9cce00006332000050e6ffffaf1a00006332;
    assign coff[418 ] = 256'h000024c8ffff856600007a9a000024c8ffffdb3800007a9affff8566ffffdb38;
    assign coff[419 ] = 256'hffff8f4d00003cafffffc351ffff8f4d000070b3ffffc35100003caf000070b3;
    assign coff[420 ] = 256'h000062b2ffffae7f00005181000062b2ffff9d4e00005181ffffae7fffff9d4e;
    assign coff[421 ] = 256'hffff8094fffff3d800000c28ffff809400007f6c00000c28fffff3d800007f6c;
    assign coff[422 ] = 256'hffffda78ffff85a000007a60ffffda780000258800007a60ffff85a000002588;
    assign coff[423 ] = 256'hffffc40200007112ffff8eeeffffc40200003bfeffff8eee0000711200003bfe;
    assign coff[424 ] = 256'h0000761bffffcea7000031590000761bffff89e500003159ffffcea7ffff89e5;
    assign coff[425 ] = 256'hffff8998ffffcf610000309fffff8998000076680000309fffffcf6100007668;
    assign coff[426 ] = 256'hffffff9bffff800100007fffffffff9b0000006500007fffffff800100000065;
    assign coff[427 ] = 256'hffffa5c500005ac9ffffa537ffffa5c500005a3bffffa53700005ac900005a3b;
    assign coff[428 ] = 256'h000046c9ffff955b00006aa5000046c9ffffb93700006aa5ffff955bffffb937;
    assign coff[429 ] = 256'hffff82890000195bffffe6a5ffff828900007d77ffffe6a50000195b00007d77;
    assign coff[430 ] = 256'hffffb890ffff95ca00006a36ffffb8900000477000006a36ffff95ca00004770;
    assign coff[431 ] = 256'hffffe76a00007d9effff8262ffffe76a00001896ffff826200007d9e00001896;
    assign coff[432 ] = 256'h00007c11ffffe08500001f7b00007c11ffff83ef00001f7bffffe085ffff83ef;
    assign coff[433 ] = 256'hffff9202ffffbe8800004178ffff920200006dfe00004178ffffbe8800006dfe;
    assign coff[434 ] = 256'h00001265ffff815400007eac00001265ffffed9b00007eacffff8154ffffed9b;
    assign coff[435 ] = 256'hffff996d00004c91ffffb36fffff996d00006693ffffb36f00004c9100006693;
    assign coff[436 ] = 256'h000055abffffa0e500005f1b000055abffffaa5500005f1bffffa0e5ffffaa55;
    assign coff[437 ] = 256'hffff802d000006acfffff954ffff802d00007fd3fffff954000006ac00007fd3;
    assign coff[438 ] = 256'hffffc8ebffff8c750000738bffffc8eb000037150000738bffff8c7500003715;
    assign coff[439 ] = 256'hffffd53f000078a6ffff875affffd53f00002ac1ffff875a000078a600002ac1;
    assign coff[440 ] = 256'h00006d96ffffbddc0000422400006d96ffff926a00004224ffffbddcffff926a;
    assign coff[441 ] = 256'hffff83beffffe14800001eb8ffff83be00007c4200001eb8ffffe14800007c42;
    assign coff[442 ] = 256'hffffecd5ffff817200007e8effffecd50000132b00007e8effff81720000132b;
    assign coff[443 ] = 256'hffffb4110000670bffff98f5ffffb41100004befffff98f50000670b00004bef;
    assign coff[444 ] = 256'h0000365fffff8c1f000073e10000365fffffc9a1000073e1ffff8c1fffffc9a1;
    assign coff[445 ] = 256'hffff879d00002b7effffd482ffff879d00007863ffffd48200002b7e00007863;
    assign coff[446 ] = 256'hffffa9c0ffffa16c00005e94ffffa9c00000564000005e94ffffa16c00005640;
    assign coff[447 ] = 256'hfffffa1d00007fddffff8023fffffa1d000005e3ffff802300007fdd000005e3;
    assign coff[448 ] = 256'h00007fbcfffff7c20000083e00007fbcffff80440000083efffff7c2ffff8044;
    assign coff[449 ] = 256'hffff9fdaffffab810000547fffff9fda000060260000547fffffab8100006026;
    assign coff[450 ] = 256'h00002945ffff86d60000792a00002945ffffd6bb0000792affff86d6ffffd6bb;
    assign coff[451 ] = 256'hffff8d240000387fffffc781ffff8d24000072dcffffc7810000387f000072dc;
    assign coff[452 ] = 256'h000065a1ffffb22f00004dd1000065a1ffff9a5f00004dd1ffffb22fffff9a5f;
    assign coff[453 ] = 256'hffff811dffffef2a000010d6ffff811d00007ee3000010d6ffffef2a00007ee3;
    assign coff[454 ] = 256'hffffdeffffff845400007bacffffdeff0000210100007bacffff845400002101;
    assign coff[455 ] = 256'hffffbfe300006ec9ffff9137ffffbfe30000401dffff913700006ec90000401d;
    assign coff[456 ] = 256'h000077d8ffffd30900002cf7000077d8ffff882800002cf7ffffd309ffff8828;
    assign coff[457 ] = 256'hffff8b77ffffcb0e000034f2ffff8b7700007489000034f2ffffcb0e00007489;
    assign coff[458 ] = 256'h00000452ffff801300007fed00000452fffffbae00007fedffff8013fffffbae;
    assign coff[459 ] = 256'hffffa27d00005767ffffa899ffffa27d00005d83ffffa8990000576700005d83;
    assign coff[460 ] = 256'h00004aaaffff9808000067f800004aaaffffb556000067f8ffff9808ffffb556;
    assign coff[461 ] = 256'hffff81b0000014b9ffffeb47ffff81b000007e50ffffeb47000014b900007e50;
    assign coff[462 ] = 256'hffffbc85ffff933c00006cc4ffffbc850000437b00006cc4ffff933c0000437b;
    assign coff[463 ] = 256'hffffe2cf00007ca0ffff8360ffffe2cf00001d31ffff836000007ca000001d31;
    assign coff[464 ] = 256'h00007d25ffffe51b00001ae500007d25ffff82db00001ae5ffffe51bffff82db;
    assign coff[465 ] = 256'hffff947effffba8700004579ffff947e00006b8200004579ffffba8700006b82;
    assign coff[466 ] = 256'h0000170bffff821700007de90000170bffffe8f500007de9ffff8217ffffe8f5;
    assign coff[467 ] = 256'hffff96ad000048bdffffb743ffff96ad00006953ffffb743000048bd00006953;
    assign coff[468 ] = 256'h0000591cffffa41d00005be30000591cffffa6e400005be3ffffa41dffffa6e4;
    assign coff[469 ] = 256'hffff8004000001f7fffffe09ffff800400007ffcfffffe09000001f700007ffc;
    assign coff[470 ] = 256'hffffcd35ffff8a820000757effffcd35000032cb0000757effff8a82000032cb;
    assign coff[471 ] = 256'hffffd0d6000076feffff8902ffffd0d600002f2affff8902000076fe00002f2a;
    assign coff[472 ] = 256'h00006ff2ffffc1f000003e1000006ff2ffff900e00003e10ffffc1f0ffff900e;
    assign coff[473 ] = 256'hffff84f5ffffdcba00002346ffff84f500007b0b00002346ffffdcba00007b0b;
    assign coff[474 ] = 256'hfffff180ffff80d300007f2dfffff18000000e8000007f2dffff80d300000e80;
    assign coff[475 ] = 256'hffffb0530000642effff9bd2ffffb05300004fadffff9bd20000642e00004fad;
    assign coff[476 ] = 256'h00003a9affff8e34000071cc00003a9affffc566000071ccffff8e34ffffc566;
    assign coff[477 ] = 256'hffff861900002708ffffd8f8ffff8619000079e7ffffd8f800002708000079e7;
    assign coff[478 ] = 256'hffffad4affff9e50000061b0ffffad4a000052b6000061b0ffff9e50000052b6;
    assign coff[479 ] = 256'hfffff56900007f90ffff8070fffff56900000a97ffff807000007f9000000a97;
    assign coff[480 ] = 256'h00007ec8ffffee620000119e00007ec8ffff81380000119effffee62ffff8138;
    assign coff[481 ] = 256'hffff99e5ffffb2cf00004d31ffff99e50000661b00004d31ffffb2cf0000661b;
    assign coff[482 ] = 256'h0000203effff842100007bdf0000203effffdfc200007bdfffff8421ffffdfc2;
    assign coff[483 ] = 256'hffff919c000040cbffffbf35ffff919c00006e64ffffbf35000040cb00006e64;
    assign coff[484 ] = 256'h00005fa1ffffaaeb0000551500005fa1ffffa05f00005515ffffaaebffffa05f;
    assign coff[485 ] = 256'hffff8038fffff88b00000775ffff803800007fc800000775fffff88b00007fc8;
    assign coff[486 ] = 256'hffffd5fdffff8717000078e9ffffd5fd00002a03000078e9ffff871700002a03;
    assign coff[487 ] = 256'hffffc83600007334ffff8cccffffc836000037caffff8ccc00007334000037ca;
    assign coff[488 ] = 256'h00007436ffffca57000035a900007436ffff8bca000035a9ffffca57ffff8bca;
    assign coff[489 ] = 256'hffff87e2ffffd3c500002c3bffff87e20000781e00002c3bffffd3c50000781e;
    assign coff[490 ] = 256'hfffffae5ffff801a00007fe6fffffae50000051b00007fe6ffff801a0000051b;
    assign coff[491 ] = 256'hffffa92c00005e0cffffa1f4ffffa92c000056d4ffffa1f400005e0c000056d4;
    assign coff[492 ] = 256'h000042d0ffff92d200006d2e000042d0ffffbd3000006d2effff92d2ffffbd30;
    assign coff[493 ] = 256'hffff838e00001df5ffffe20bffff838e00007c72ffffe20b00001df500007c72;
    assign coff[494 ] = 256'hffffb4b3ffff987e00006782ffffb4b300004b4d00006782ffff987e00004b4d;
    assign coff[495 ] = 256'hffffec0e00007e70ffff8190ffffec0e000013f2ffff819000007e70000013f2;
    assign coff[496 ] = 256'h00007ad3ffffdbf90000240700007ad3ffff852d00002407ffffdbf9ffff852d;
    assign coff[497 ] = 256'hffff8fadffffc2a000003d60ffff8fad0000705300003d60ffffc2a000007053;
    assign coff[498 ] = 256'h00000db8ffff80bd00007f4300000db8fffff24800007f43ffff80bdfffff248;
    assign coff[499 ] = 256'hffff9c500000504affffafb6ffff9c50000063b0ffffafb60000504a000063b0;
    assign coff[500 ] = 256'h0000521cffff9dce000062320000521cffffade400006232ffff9dceffffade4;
    assign coff[501 ] = 256'hffff808200000b60fffff4a0ffff808200007f7efffff4a000000b6000007f7e;
    assign coff[502 ] = 256'hffffc4b4ffff8e9000007170ffffc4b400003b4c00007170ffff8e9000003b4c;
    assign coff[503 ] = 256'hffffd9b800007a24ffff85dcffffd9b800002648ffff85dc00007a2400002648;
    assign coff[504 ] = 256'h00006b14ffffb9df0000462100006b14ffff94ec00004621ffffb9dfffff94ec;
    assign coff[505 ] = 256'hffff82b2ffffe5e000001a20ffff82b200007d4e00001a20ffffe5e000007d4e;
    assign coff[506 ] = 256'hffffe82fffff823c00007dc4ffffe82f000017d100007dc4ffff823c000017d1;
    assign coff[507 ] = 256'hffffb7e9000069c5ffff963bffffb7e900004817ffff963b000069c500004817;
    assign coff[508 ] = 256'h00003212ffff8a33000075cd00003212ffffcdee000075cdffff8a33ffffcdee;
    assign coff[509 ] = 256'hffff894c00002fe5ffffd01bffff894c000076b4ffffd01b00002fe5000076b4;
    assign coff[510 ] = 256'hffffa654ffffa4a900005b57ffffa654000059ac00005b57ffffa4a9000059ac;
    assign coff[511 ] = 256'hfffffed200007fffffff8001fffffed20000012effff800100007fff0000012e;
    assign coff[512 ] = 256'h00007fffffffff690000009700007fffffff800100000097ffffff69ffff8001;
    assign coff[513 ] = 256'hffffa513ffffa5e800005a18ffffa51300005aed00005a18ffffa5e800005aed;
    assign coff[514 ] = 256'h00003070ffff89850000767b00003070ffffcf900000767bffff8985ffffcf90;
    assign coff[515 ] = 256'hffff89f800003187ffffce79ffff89f800007608ffffce790000318700007608;
    assign coff[516 ] = 256'h00006a1affffb8660000479a00006a1affff95e60000479affffb866ffff95e6;
    assign coff[517 ] = 256'hffff8259ffffe79b00001865ffff825900007da700001865ffffe79b00007da7;
    assign coff[518 ] = 256'hffffe673ffff829300007d6dffffe6730000198d00007d6dffff82930000198d;
    assign coff[519 ] = 256'hffffb96100006ac1ffff953fffffb9610000469fffff953f00006ac10000469f;
    assign coff[520 ] = 256'h00007a51ffffda48000025b800007a51ffff85af000025b8ffffda48ffff85af;
    assign coff[521 ] = 256'hffff8ed6ffffc42e00003bd2ffff8ed60000712a00003bd2ffffc42e0000712a;
    assign coff[522 ] = 256'h00000bf6ffff808f00007f7100000bf6fffff40a00007f71ffff808ffffff40a;
    assign coff[523 ] = 256'hffff9d6e000051a8ffffae58ffff9d6e00006292ffffae58000051a800006292;
    assign coff[524 ] = 256'h000050bfffff9caf00006351000050bfffffaf4100006351ffff9cafffffaf41;
    assign coff[525 ] = 256'hffff80ad00000d22fffff2deffff80ad00007f53fffff2de00000d2200007f53;
    assign coff[526 ] = 256'hffffc324ffff8f650000709bffffc32400003cdc0000709bffff8f6500003cdc;
    assign coff[527 ] = 256'hffffdb6800007aa8ffff8558ffffdb6800002498ffff855800007aa800002498;
    assign coff[528 ] = 256'h00007e87ffffeca30000135d00007e87ffff81790000135dffffeca3ffff8179;
    assign coff[529 ] = 256'hffff98d7ffffb43900004bc7ffff98d70000672900004bc7ffffb43900006729;
    assign coff[530 ] = 256'h00001e88ffff83b200007c4e00001e88ffffe17800007c4effff83b2ffffe178;
    assign coff[531 ] = 256'hffff92840000424fffffbdb1ffff928400006d7cffffbdb10000424f00006d7c;
    assign coff[532 ] = 256'h00005e72ffffa99b0000566500005e72ffffa18e00005665ffffa99bffffa18e;
    assign coff[533 ] = 256'hffff8020fffffa4f000005b1ffff802000007fe0000005b1fffffa4f00007fe0;
    assign coff[534 ] = 256'hffffd453ffff87af00007851ffffd45300002bad00007851ffff87af00002bad;
    assign coff[535 ] = 256'hffffc9ce000073f6ffff8c0affffc9ce00003632ffff8c0a000073f600003632;
    assign coff[536 ] = 256'h00007375ffffc8be0000374200007375ffff8c8b00003742ffffc8beffff8c8b;
    assign coff[537 ] = 256'hffff8749ffffd56f00002a91ffff8749000078b700002a91ffffd56f000078b7;
    assign coff[538 ] = 256'hfffff922ffff802f00007fd1fffff922000006de00007fd1ffff802f000006de;
    assign coff[539 ] = 256'hffffaa7a00005f3cffffa0c4ffffaa7a00005586ffffa0c400005f3c00005586;
    assign coff[540 ] = 256'h0000414dffff91e900006e170000414dffffbeb300006e17ffff91e9ffffbeb3;
    assign coff[541 ] = 256'hffff83fb00001facffffe054ffff83fb00007c05ffffe05400001fac00007c05;
    assign coff[542 ] = 256'hffffb347ffff998b00006675ffffb34700004cb900006675ffff998b00004cb9;
    assign coff[543 ] = 256'hffffedcd00007eb3ffff814dffffedcd00001233ffff814d00007eb300001233;
    assign coff[544 ] = 256'h00007f9cfffff5ff00000a0100007f9cffff806400000a01fffff5ffffff8064;
    assign coff[545 ] = 256'hffff9eb2ffffacd700005329ffff9eb20000614e00005329ffffacd70000614e;
    assign coff[546 ] = 256'h00002797ffff8647000079b900002797ffffd869000079b9ffff8647ffffd869;
    assign coff[547 ] = 256'hffff8def00003a13ffffc5edffff8def00007211ffffc5ed00003a1300007211;
    assign coff[548 ] = 256'h0000648bffffb0c900004f370000648bffff9b7500004f37ffffb0c9ffff9b75;
    assign coff[549 ] = 256'hffff80e4fffff0eb00000f15ffff80e400007f1c00000f15fffff0eb00007f1c;
    assign coff[550 ] = 256'hffffdd4bffff84cc00007b34ffffdd4b000022b500007b34ffff84cc000022b5;
    assign coff[551 ] = 256'hffffc16c00006fa9ffff9057ffffc16c00003e94ffff905700006fa900003e94;
    assign coff[552 ] = 256'h00007736ffffd16200002e9e00007736ffff88ca00002e9effffd162ffff88ca;
    assign coff[553 ] = 256'hffff8abeffffccab00003355ffff8abe0000754200003355ffffccab00007542;
    assign coff[554 ] = 256'h0000028dffff800700007ff90000028dfffffd7300007ff9ffff8007fffffd73;
    assign coff[555 ] = 256'hffffa3b4000058b0ffffa750ffffa3b400005c4cffffa750000058b000005c4c;
    assign coff[556 ] = 256'h00004939ffff9703000068fd00004939ffffb6c7000068fdffff9703ffffb6c7;
    assign coff[557 ] = 256'hffff81fd00001677ffffe989ffff81fd00007e03ffffe9890000167700007e03;
    assign coff[558 ] = 256'hffffbb06ffff942d00006bd3ffffbb06000044fa00006bd3ffff942d000044fa;
    assign coff[559 ] = 256'hffffe48800007d05ffff82fbffffe48800001b78ffff82fb00007d0500001b78;
    assign coff[560 ] = 256'h00007cc2ffffe36100001c9f00007cc2ffff833e00001c9fffffe361ffff833e;
    assign coff[561 ] = 256'hffff938bffffbc05000043fbffff938b00006c75000043fbffffbc0500006c75;
    assign coff[562 ] = 256'h0000154dffff81c900007e370000154dffffeab300007e37ffff81c9ffffeab3;
    assign coff[563 ] = 256'hffff97b000004a2fffffb5d1ffff97b000006850ffffb5d100004a2f00006850;
    assign coff[564 ] = 256'h000057d5ffffa2e400005d1c000057d5ffffa82b00005d1cffffa2e4ffffa82b;
    assign coff[565 ] = 256'hffff800e000003bbfffffc45ffff800e00007ff2fffffc45000003bb00007ff2;
    assign coff[566 ] = 256'hffffcb97ffff8b39000074c7ffffcb9700003469000074c7ffff8b3900003469;
    assign coff[567 ] = 256'hffffd27c000077a2ffff885effffd27c00002d84ffff885e000077a200002d84;
    assign coff[568 ] = 256'h00006f14ffffc06600003f9a00006f14ffff90ec00003f9affffc066ffff90ec;
    assign coff[569 ] = 256'hffff847bffffde6e00002192ffff847b00007b8500002192ffffde6e00007b85;
    assign coff[570 ] = 256'hffffefbfffff810900007ef7ffffefbf0000104100007ef7ffff810900001041;
    assign coff[571 ] = 256'hffffb1b700006545ffff9abbffffb1b700004e49ffff9abb0000654500004e49;
    assign coff[572 ] = 256'h00003906ffff8d670000729900003906ffffc6fa00007299ffff8d67ffffc6fa;
    assign coff[573 ] = 256'hffff86a5000028b6ffffd74affff86a50000795bffffd74a000028b60000795b;
    assign coff[574 ] = 256'hffffabf3ffff9f7700006089ffffabf30000540d00006089ffff9f770000540d;
    assign coff[575 ] = 256'hfffff72c00007fb2ffff804efffff72c000008d4ffff804e00007fb2000008d4;
    assign coff[576 ] = 256'h00007fe4fffffab30000054d00007fe4ffff801c0000054dfffffab3ffff801c;
    assign coff[577 ] = 256'hffffa1d2ffffa951000056afffffa1d200005e2e000056afffffa95100005e2e;
    assign coff[578 ] = 256'h00002c0cffff87d10000782f00002c0cffffd3f40000782fffff87d1ffffd3f4;
    assign coff[579 ] = 256'hffff8bdf000035d7ffffca29ffff8bdf00007421ffffca29000035d700007421;
    assign coff[580 ] = 256'h00006764ffffb48b00004b7500006764ffff989c00004b75ffffb48bffff989c;
    assign coff[581 ] = 256'hffff8188ffffec3f000013c1ffff818800007e78000013c1ffffec3f00007e78;
    assign coff[582 ] = 256'hffffe1daffff839a00007c66ffffe1da00001e2600007c66ffff839a00001e26;
    assign coff[583 ] = 256'hffffbd5b00006d48ffff92b8ffffbd5b000042a5ffff92b800006d48000042a5;
    assign coff[584 ] = 256'h000078d8ffffd5ce00002a32000078d8ffff872800002a32ffffd5ceffff8728;
    assign coff[585 ] = 256'hffff8cb6ffffc8630000379dffff8cb60000734a0000379dffffc8630000734a;
    assign coff[586 ] = 256'h00000743ffff803500007fcb00000743fffff8bd00007fcbffff8035fffff8bd;
    assign coff[587 ] = 256'hffffa0800000553bffffaac5ffffa08000005f80ffffaac50000553b00005f80;
    assign coff[588 ] = 256'h00004d09ffff99c70000663900004d09ffffb2f700006639ffff99c7ffffb2f7;
    assign coff[589 ] = 256'hffff813f000011cfffffee31ffff813f00007ec1ffffee31000011cf00007ec1;
    assign coff[590 ] = 256'hffffbf0affff91b600006e4affffbf0a000040f600006e4affff91b6000040f6;
    assign coff[591 ] = 256'hffffdff200007becffff8414ffffdff20000200effff841400007bec0000200e;
    assign coff[592 ] = 256'h00007dbaffffe7fe0000180200007dbaffff824600001802ffffe7feffff8246;
    assign coff[593 ] = 256'hffff961fffffb813000047edffff961f000069e1000047edffffb813000069e1;
    assign coff[594 ] = 256'h000019efffff82a800007d58000019efffffe61100007d58ffff82a8ffffe611;
    assign coff[595 ] = 256'hffff95080000464bffffb9b5ffff950800006af8ffffb9b50000464b00006af8;
    assign coff[596 ] = 256'h00005b34ffffa630000059d000005b34ffffa4cc000059d0ffffa630ffffa4cc;
    assign coff[597 ] = 256'hffff8001ffffff05000000fbffff800100007fff000000fbffffff0500007fff;
    assign coff[598 ] = 256'hffffcfedffff895f000076a1ffffcfed00003013000076a1ffff895f00003013;
    assign coff[599 ] = 256'hffffce1c000075e1ffff8a1fffffce1c000031e4ffff8a1f000075e1000031e4;
    assign coff[600 ] = 256'h00007158ffffc48700003b7900007158ffff8ea800003b79ffffc487ffff8ea8;
    assign coff[601 ] = 256'hffff85cdffffd9e800002618ffff85cd00007a3300002618ffffd9e800007a33;
    assign coff[602 ] = 256'hfffff46effff808600007f7afffff46e00000b9200007f7affff808600000b92;
    assign coff[603 ] = 256'hffffae0b00006252ffff9daeffffae0b000051f5ffff9dae00006252000051f5;
    assign coff[604 ] = 256'h00003d34ffff8f950000706b00003d34ffffc2cc0000706bffff8f95ffffc2cc;
    assign coff[605 ] = 256'hffff853b00002437ffffdbc9ffff853b00007ac5ffffdbc90000243700007ac5;
    assign coff[606 ] = 256'hffffaf8fffff9c6f00006391ffffaf8f0000507100006391ffff9c6f00005071;
    assign coff[607 ] = 256'hfffff27a00007f49ffff80b7fffff27a00000d86ffff80b700007f4900000d86;
    assign coff[608 ] = 256'h00007f27fffff14e00000eb200007f27ffff80d900000eb2fffff14effff80d9;
    assign coff[609 ] = 256'hffff9bb3ffffb07b00004f85ffff9bb30000644d00004f85ffffb07b0000644d;
    assign coff[610 ] = 256'h00002316ffff84e700007b1900002316ffffdcea00007b19ffff84e7ffffdcea;
    assign coff[611 ] = 256'hffff902600003e3cffffc1c4ffff902600006fdaffffc1c400003e3c00006fda;
    assign coff[612 ] = 256'h00006190ffffad24000052dc00006190ffff9e70000052dcffffad24ffff9e70;
    assign coff[613 ] = 256'hffff806cfffff59b00000a65ffff806c00007f9400000a65fffff59b00007f94;
    assign coff[614 ] = 256'hffffd8c8ffff8628000079d8ffffd8c800002738000079d8ffff862800002738;
    assign coff[615 ] = 256'hffffc593000071e3ffff8e1dffffc59300003a6dffff8e1d000071e300003a6d;
    assign coff[616 ] = 256'h0000756affffcd07000032f90000756affff8a96000032f9ffffcd07ffff8a96;
    assign coff[617 ] = 256'hffff88efffffd10500002efbffff88ef0000771100002efbffffd10500007711;
    assign coff[618 ] = 256'hfffffdd7ffff800500007ffbfffffdd70000022900007ffbffff800500000229;
    assign coff[619 ] = 256'hffffa70800005c06ffffa3faffffa708000058f8ffffa3fa00005c06000058f8;
    assign coff[620 ] = 256'h0000454fffff946300006b9d0000454fffffbab100006b9dffff9463ffffbab1;
    assign coff[621 ] = 256'hffff82e600001b16ffffe4eaffff82e600007d1affffe4ea00001b1600007d1a;
    assign coff[622 ] = 256'hffffb71affff96c900006937ffffb71a000048e600006937ffff96c9000048e6;
    assign coff[623 ] = 256'hffffe92600007df2ffff820effffe926000016daffff820e00007df2000016da;
    assign coff[624 ] = 256'h00007b9fffffdecf0000213100007b9fffff846100002131ffffdecfffff8461;
    assign coff[625 ] = 256'hffff911effffc00f00003ff1ffff911e00006ee200003ff1ffffc00f00006ee2;
    assign coff[626 ] = 256'h000010a4ffff811600007eea000010a4ffffef5c00007eeaffff8116ffffef5c;
    assign coff[627 ] = 256'hffff9a7e00004df9ffffb207ffff9a7e00006582ffffb20700004df900006582;
    assign coff[628 ] = 256'h00005459ffff9fb90000604700005459ffffaba700006047ffff9fb9ffffaba7;
    assign coff[629 ] = 256'hffff804700000870fffff790ffff804700007fb9fffff7900000087000007fb9;
    assign coff[630 ] = 256'hffffc754ffff8d3b000072c5ffffc754000038ac000072c5ffff8d3b000038ac;
    assign coff[631 ] = 256'hffffd6eb0000793affff86c6ffffd6eb00002915ffff86c60000793a00002915;
    assign coff[632 ] = 256'h00006caaffffbc5a000043a600006caaffff9356000043a6ffffbc5affff9356;
    assign coff[633 ] = 256'hffff8354ffffe2ff00001d01ffff835400007cac00001d01ffffe2ff00007cac;
    assign coff[634 ] = 256'hffffeb16ffff81b800007e48ffffeb16000014ea00007e48ffff81b8000014ea;
    assign coff[635 ] = 256'hffffb57f00006815ffff97ebffffb57f00004a81ffff97eb0000681500004a81;
    assign coff[636 ] = 256'h000034c4ffff8b620000749e000034c4ffffcb3c0000749effff8b62ffffcb3c;
    assign coff[637 ] = 256'hffff883a00002d26ffffd2daffff883a000077c6ffffd2da00002d26000077c6;
    assign coff[638 ] = 256'hffffa874ffffa29f00005d61ffffa8740000578c00005d61ffffa29f0000578c;
    assign coff[639 ] = 256'hfffffbe100007fefffff8011fffffbe10000041fffff801100007fef0000041f;
    assign coff[640 ] = 256'h00007ff7fffffd0e000002f200007ff7ffff8009000002f2fffffd0effff8009;
    assign coff[641 ] = 256'hffffa36fffffa79900005867ffffa36f00005c9100005867ffffa79900005c91;
    assign coff[642 ] = 256'h00002e40ffff88a60000775a00002e40ffffd1c00000775affff88a6ffffd1c0;
    assign coff[643 ] = 256'hffff8ae7000033b1ffffcc4fffff8ae700007519ffffcc4f000033b100007519;
    assign coff[644 ] = 256'h000068c4ffffb6750000498b000068c4ffff973c0000498bffffb675ffff973c;
    assign coff[645 ] = 256'hffff81ebffffe9ec00001614ffff81eb00007e1500001614ffffe9ec00007e15;
    assign coff[646 ] = 256'hffffe426ffff831100007cefffffe42600001bda00007cefffff831100001bda;
    assign coff[647 ] = 256'hffffbb5b00006c09ffff93f7ffffbb5b000044a5ffff93f700006c09000044a5;
    assign coff[648 ] = 256'h0000799affffd809000027f70000799affff8666000027f7ffffd809ffff8666;
    assign coff[649 ] = 256'hffff8dc1ffffc646000039baffff8dc10000723f000039baffffc6460000723f;
    assign coff[650 ] = 256'h0000099dffff805d00007fa30000099dfffff66300007fa3ffff805dfffff663;
    assign coff[651 ] = 256'hffff9ef300005375ffffac8bffff9ef30000610dffffac8b000053750000610d;
    assign coff[652 ] = 256'h00004ee8ffff9b36000064ca00004ee8ffffb118000064caffff9b36ffffb118;
    assign coff[653 ] = 256'hffff80f000000f79fffff087ffff80f000007f10fffff08700000f7900007f10;
    assign coff[654 ] = 256'hffffc114ffff908800006f78ffffc11400003eec00006f78ffff908800003eec;
    assign coff[655 ] = 256'hffffddac00007b50ffff84b0ffffddac00002254ffff84b000007b5000002254;
    assign coff[656 ] = 256'h00007e26ffffea4f000015b100007e26ffff81da000015b1ffffea4fffff81da;
    assign coff[657 ] = 256'hffff9776ffffb623000049ddffff97760000688a000049ddffffb6230000688a;
    assign coff[658 ] = 256'h00001c3dffff832700007cd900001c3dffffe3c300007cd9ffff8327ffffe3c3;
    assign coff[659 ] = 256'hffff93c100004450ffffbbb0ffff93c100006c3fffffbbb00000445000006c3f;
    assign coff[660 ] = 256'h00005cd7ffffa7e20000581e00005cd7ffffa3290000581effffa7e2ffffa329;
    assign coff[661 ] = 256'hffff800bfffffcaa00000356ffff800b00007ff500000356fffffcaa00007ff5;
    assign coff[662 ] = 256'hffffd21effff88820000777effffd21e00002de20000777effff888200002de2;
    assign coff[663 ] = 256'hffffcbf3000074f0ffff8b10ffffcbf30000340dffff8b10000074f00000340d;
    assign coff[664 ] = 256'h0000726cffffc6a0000039600000726cffff8d9400003960ffffc6a0ffff8d94;
    assign coff[665 ] = 256'hffff8686ffffd7aa00002856ffff86860000797a00002856ffffd7aa0000797a;
    assign coff[666 ] = 256'hfffff6c8ffff805500007fabfffff6c80000093800007fabffff805500000938;
    assign coff[667 ] = 256'hffffac3f000060cbffff9f35ffffac3f000053c1ffff9f35000060cb000053c1;
    assign coff[668 ] = 256'h00003f43ffff90ba00006f4600003f43ffffc0bd00006f46ffff90baffffc0bd;
    assign coff[669 ] = 256'hffff8496000021f3ffffde0dffff849600007b6affffde0d000021f300007b6a;
    assign coff[670 ] = 256'hffffb168ffff9af900006507ffffb16800004e9800006507ffff9af900004e98;
    assign coff[671 ] = 256'hfffff02300007f03ffff80fdfffff02300000fddffff80fd00007f0300000fdd;
    assign coff[672 ] = 256'h00007f67fffff3a600000c5a00007f67ffff809900000c5afffff3a6ffff8099;
    assign coff[673 ] = 256'hffff9d2effffaea50000515bffff9d2e000062d20000515bffffaea5000062d2;
    assign coff[674 ] = 256'h00002558ffff859200007a6e00002558ffffdaa800007a6effff8592ffffdaa8;
    assign coff[675 ] = 256'hffff8f0600003c2affffc3d6ffff8f06000070faffffc3d600003c2a000070fa;
    assign coff[676 ] = 256'h00006312ffffaef30000510d00006312ffff9cee0000510dffffaef3ffff9cee;
    assign coff[677 ] = 256'hffff80a3fffff34200000cbeffff80a300007f5d00000cbefffff34200007f5d;
    assign coff[678 ] = 256'hffffdb08ffff857400007a8cffffdb08000024f800007a8cffff8574000024f8;
    assign coff[679 ] = 256'hffffc37d000070cbffff8f35ffffc37d00003c83ffff8f35000070cb00003c83;
    assign coff[680 ] = 256'h00007655ffffcf33000030cd00007655ffff89ab000030cdffffcf33ffff89ab;
    assign coff[681 ] = 256'hffff89d2ffffced60000312affff89d20000762e0000312affffced60000762e;
    assign coff[682 ] = 256'h00000032ffff800100007fff00000032ffffffce00007fffffff8001ffffffce;
    assign coff[683 ] = 256'hffffa55a00005a5fffffa5a1ffffa55a00005aa6ffffa5a100005a5f00005aa6;
    assign coff[684 ] = 256'h00004747ffff95ae00006a5200004747ffffb8b900006a52ffff95aeffffb8b9;
    assign coff[685 ] = 256'hffff826c000018c7ffffe739ffff826c00007d94ffffe739000018c700007d94;
    assign coff[686 ] = 256'hffffb90dffff957700006a89ffffb90d000046f300006a89ffff9577000046f3;
    assign coff[687 ] = 256'hffffe6d600007d81ffff827fffffe6d60000192affff827f00007d810000192a;
    assign coff[688 ] = 256'h00007c36ffffe11700001ee900007c36ffff83ca00001ee9ffffe117ffff83ca;
    assign coff[689 ] = 256'hffff9250ffffbe07000041f9ffff925000006db0000041f9ffffbe0700006db0;
    assign coff[690 ] = 256'h000012faffff816a00007e96000012faffffed0600007e96ffff816affffed06;
    assign coff[691 ] = 256'hffff991300004c17ffffb3e9ffff9913000066edffffb3e900004c17000066ed;
    assign coff[692 ] = 256'h0000561bffffa14a00005eb60000561bffffa9e500005eb6ffffa14affffa9e5;
    assign coff[693 ] = 256'hffff802500000616fffff9eaffff802500007fdbfffff9ea0000061600007fdb;
    assign coff[694 ] = 256'hffffc973ffff8c35000073cbffffc9730000368d000073cbffff8c350000368d;
    assign coff[695 ] = 256'hffffd4b100007874ffff878cffffd4b100002b4fffff878c0000787400002b4f;
    assign coff[696 ] = 256'h00006de4ffffbe5d000041a300006de4ffff921c000041a3ffffbe5dffff921c;
    assign coff[697 ] = 256'hffff83e2ffffe0b500001f4bffff83e200007c1e00001f4bffffe0b500007c1e;
    assign coff[698 ] = 256'hffffed6affff815b00007ea5ffffed6a0000129600007ea5ffff815b00001296;
    assign coff[699 ] = 256'hffffb398000066b2ffff994effffb39800004c68ffff994e000066b200004c68;
    assign coff[700 ] = 256'h000036e8ffff8c60000073a0000036e8ffffc918000073a0ffff8c60ffffc918;
    assign coff[701 ] = 256'hffff876b00002af0ffffd510ffff876b00007895ffffd51000002af000007895;
    assign coff[702 ] = 256'hffffaa30ffffa10700005ef9ffffaa30000055d000005ef9ffffa107000055d0;
    assign coff[703 ] = 256'hfffff98600007fd6ffff802afffff9860000067affff802a00007fd60000067a;
    assign coff[704 ] = 256'h00007fc5fffff859000007a700007fc5ffff803b000007a7fffff859ffff803b;
    assign coff[705 ] = 256'hffffa03effffab10000054f0ffffa03e00005fc2000054f0ffffab1000005fc2;
    assign coff[706 ] = 256'h000029d3ffff8707000078f9000029d3ffffd62d000078f9ffff8707ffffd62d;
    assign coff[707 ] = 256'hffff8ce2000037f7ffffc809ffff8ce20000731effffc809000037f70000731e;
    assign coff[708 ] = 256'h000065fcffffb2a700004d59000065fcffff9a0400004d59ffffb2a7ffff9a04;
    assign coff[709 ] = 256'hffff8131ffffee940000116cffff813100007ecf0000116cffffee9400007ecf;
    assign coff[710 ] = 256'hffffdf91ffff842d00007bd3ffffdf910000206f00007bd3ffff842d0000206f;
    assign coff[711 ] = 256'hffffbf6100006e7dffff9183ffffbf610000409fffff918300006e7d0000409f;
    assign coff[712 ] = 256'h0000780cffffd39600002c6a0000780cffff87f400002c6affffd396ffff87f4;
    assign coff[713 ] = 256'hffff8bb5ffffca850000357bffff8bb50000744b0000357bffffca850000744b;
    assign coff[714 ] = 256'h000004e8ffff801800007fe8000004e8fffffb1800007fe8ffff8018fffffb18;
    assign coff[715 ] = 256'hffffa216000056f9ffffa907ffffa21600005deaffffa907000056f900005dea;
    assign coff[716 ] = 256'h00004b24ffff9860000067a000004b24ffffb4dc000067a0ffff9860ffffb4dc;
    assign coff[717 ] = 256'hffff819800001424ffffebdcffff819800007e68ffffebdc0000142400007e68;
    assign coff[718 ] = 256'hffffbd05ffff92ec00006d14ffffbd05000042fb00006d14ffff92ec000042fb;
    assign coff[719 ] = 256'hffffe23c00007c7effff8382ffffe23c00001dc4ffff838200007c7e00001dc4;
    assign coff[720 ] = 256'h00007d44ffffe5af00001a5100007d44ffff82bc00001a51ffffe5afffff82bc;
    assign coff[721 ] = 256'hffff94d0ffffba09000045f7ffff94d000006b30000045f7ffffba0900006b30;
    assign coff[722 ] = 256'h0000179fffff823300007dcd0000179fffffe86100007dcdffff8233ffffe861;
    assign coff[723 ] = 256'hffff965700004840ffffb7c0ffff9657000069a9ffffb7c000004840000069a9;
    assign coff[724 ] = 256'h00005988ffffa48600005b7a00005988ffffa67800005b7affffa486ffffa678;
    assign coff[725 ] = 256'hffff800200000160fffffea0ffff800200007ffefffffea00000016000007ffe;
    assign coff[726 ] = 256'hffffcdc0ffff8a47000075b9ffffcdc000003240000075b9ffff8a4700003240;
    assign coff[727 ] = 256'hffffd04a000076c7ffff8939ffffd04a00002fb6ffff8939000076c700002fb6;
    assign coff[728 ] = 256'h0000703bffffc27400003d8c0000703bffff8fc500003d8cffffc274ffff8fc5;
    assign coff[729 ] = 256'hffff851fffffdc29000023d7ffff851f00007ae1000023d7ffffdc2900007ae1;
    assign coff[730 ] = 256'hfffff216ffff80c200007f3efffff21600000dea00007f3effff80c200000dea;
    assign coff[731 ] = 256'hffffafdd000063d0ffff9c30ffffafdd00005023ffff9c30000063d000005023;
    assign coff[732 ] = 256'h00003b20ffff8e790000718700003b20ffffc4e000007187ffff8e79ffffc4e0;
    assign coff[733 ] = 256'hffff85eb00002678ffffd988ffff85eb00007a15ffffd9880000267800007a15;
    assign coff[734 ] = 256'hffffadbdffff9def00006211ffffadbd0000524300006211ffff9def00005243;
    assign coff[735 ] = 256'hfffff4d300007f83ffff807dfffff4d300000b2dffff807d00007f8300000b2d;
    assign coff[736 ] = 256'h00007eddffffeef80000110800007eddffff812300001108ffffeef8ffff8123;
    assign coff[737 ] = 256'hffff9a40ffffb25700004da9ffff9a40000065c000004da9ffffb257000065c0;
    assign coff[738 ] = 256'h000020d0ffff844700007bb9000020d0ffffdf3000007bb9ffff8447ffffdf30;
    assign coff[739 ] = 256'hffff915000004048ffffbfb8ffff915000006eb0ffffbfb80000404800006eb0;
    assign coff[740 ] = 256'h00006005ffffab5c000054a400006005ffff9ffb000054a4ffffab5cffff9ffb;
    assign coff[741 ] = 256'hffff8041fffff7f40000080cffff804100007fbf0000080cfffff7f400007fbf;
    assign coff[742 ] = 256'hffffd68cffff86e60000791affffd68c000029740000791affff86e600002974;
    assign coff[743 ] = 256'hffffc7ae000072f2ffff8d0effffc7ae00003852ffff8d0e000072f200003852;
    assign coff[744 ] = 256'h00007475ffffcae00000352000007475ffff8b8b00003520ffffcae0ffff8b8b;
    assign coff[745 ] = 256'hffff8817ffffd33800002cc8ffff8817000077e900002cc8ffffd338000077e9;
    assign coff[746 ] = 256'hfffffb7cffff801400007fecfffffb7c0000048400007fecffff801400000484;
    assign coff[747 ] = 256'hffffa8bd00005da5ffffa25bffffa8bd00005743ffffa25b00005da500005743;
    assign coff[748 ] = 256'h00004351ffff932100006cdf00004351ffffbcaf00006cdfffff9321ffffbcaf;
    assign coff[749 ] = 256'hffff836b00001d62ffffe29effff836b00007c95ffffe29e00001d6200007c95;
    assign coff[750 ] = 256'hffffb52dffff9826000067daffffb52d00004ad3000067daffff982600004ad3;
    assign coff[751 ] = 256'hffffeb7900007e58ffff81a8ffffeb7900001487ffff81a800007e5800001487;
    assign coff[752 ] = 256'h00007afdffffdc8a0000237600007afdffff850300002376ffffdc8affff8503;
    assign coff[753 ] = 256'hffff8ff5ffffc21c00003de4ffff8ff50000700b00003de4ffffc21c0000700b;
    assign coff[754 ] = 256'h00000e4effff80cd00007f3300000e4efffff1b200007f33ffff80cdfffff1b2;
    assign coff[755 ] = 256'hffff9bf100004fd4ffffb02cffff9bf10000640fffffb02c00004fd40000640f;
    assign coff[756 ] = 256'h00005290ffff9e2f000061d100005290ffffad70000061d1ffff9e2fffffad70;
    assign coff[757 ] = 256'hffff807500000ac9fffff537ffff807500007f8bfffff53700000ac900007f8b;
    assign coff[758 ] = 256'hffffc53affff8e4b000071b5ffffc53a00003ac6000071b5ffff8e4b00003ac6;
    assign coff[759 ] = 256'hffffd928000079f7ffff8609ffffd928000026d8ffff8609000079f7000026d8;
    assign coff[760 ] = 256'h00006b66ffffba5d000045a300006b66ffff949a000045a3ffffba5dffff949a;
    assign coff[761 ] = 256'hffff82d1ffffe54c00001ab4ffff82d100007d2f00001ab4ffffe54c00007d2f;
    assign coff[762 ] = 256'hffffe8c4ffff822000007de0ffffe8c40000173c00007de0ffff82200000173c;
    assign coff[763 ] = 256'hffffb76d00006970ffff9690ffffb76d00004893ffff96900000697000004893;
    assign coff[764 ] = 256'h0000329dffff8a6e000075920000329dffffcd6300007592ffff8a6effffcd63;
    assign coff[765 ] = 256'hffff891400002f59ffffd0a7ffff8914000076ecffffd0a700002f59000076ec;
    assign coff[766 ] = 256'hffffa6c0ffffa44000005bc0ffffa6c00000594000005bc0ffffa44000005940;
    assign coff[767 ] = 256'hfffffe3c00007ffdffff8003fffffe3c000001c4ffff800300007ffd000001c4;
    assign coff[768 ] = 256'h00007ffdfffffe3c000001c400007ffdffff8003000001c4fffffe3cffff8003;
    assign coff[769 ] = 256'hffffa440ffffa6c000005940ffffa44000005bc000005940ffffa6c000005bc0;
    assign coff[770 ] = 256'h00002f59ffff8914000076ec00002f59ffffd0a7000076ecffff8914ffffd0a7;
    assign coff[771 ] = 256'hffff8a6e0000329dffffcd63ffff8a6e00007592ffffcd630000329d00007592;
    assign coff[772 ] = 256'h00006970ffffb76d0000489300006970ffff969000004893ffffb76dffff9690;
    assign coff[773 ] = 256'hffff8220ffffe8c40000173cffff822000007de00000173cffffe8c400007de0;
    assign coff[774 ] = 256'hffffe54cffff82d100007d2fffffe54c00001ab400007d2fffff82d100001ab4;
    assign coff[775 ] = 256'hffffba5d00006b66ffff949affffba5d000045a3ffff949a00006b66000045a3;
    assign coff[776 ] = 256'h000079f7ffffd928000026d8000079f7ffff8609000026d8ffffd928ffff8609;
    assign coff[777 ] = 256'hffff8e4bffffc53a00003ac6ffff8e4b000071b500003ac6ffffc53a000071b5;
    assign coff[778 ] = 256'h00000ac9ffff807500007f8b00000ac9fffff53700007f8bffff8075fffff537;
    assign coff[779 ] = 256'hffff9e2f00005290ffffad70ffff9e2f000061d1ffffad7000005290000061d1;
    assign coff[780 ] = 256'h00004fd4ffff9bf10000640f00004fd4ffffb02c0000640fffff9bf1ffffb02c;
    assign coff[781 ] = 256'hffff80cd00000e4efffff1b2ffff80cd00007f33fffff1b200000e4e00007f33;
    assign coff[782 ] = 256'hffffc21cffff8ff50000700bffffc21c00003de40000700bffff8ff500003de4;
    assign coff[783 ] = 256'hffffdc8a00007afdffff8503ffffdc8a00002376ffff850300007afd00002376;
    assign coff[784 ] = 256'h00007e58ffffeb790000148700007e58ffff81a800001487ffffeb79ffff81a8;
    assign coff[785 ] = 256'hffff9826ffffb52d00004ad3ffff9826000067da00004ad3ffffb52d000067da;
    assign coff[786 ] = 256'h00001d62ffff836b00007c9500001d62ffffe29e00007c95ffff836bffffe29e;
    assign coff[787 ] = 256'hffff932100004351ffffbcafffff932100006cdfffffbcaf0000435100006cdf;
    assign coff[788 ] = 256'h00005da5ffffa8bd0000574300005da5ffffa25b00005743ffffa8bdffffa25b;
    assign coff[789 ] = 256'hffff8014fffffb7c00000484ffff801400007fec00000484fffffb7c00007fec;
    assign coff[790 ] = 256'hffffd338ffff8817000077e9ffffd33800002cc8000077e9ffff881700002cc8;
    assign coff[791 ] = 256'hffffcae000007475ffff8b8bffffcae000003520ffff8b8b0000747500003520;
    assign coff[792 ] = 256'h000072f2ffffc7ae00003852000072f2ffff8d0e00003852ffffc7aeffff8d0e;
    assign coff[793 ] = 256'hffff86e6ffffd68c00002974ffff86e60000791a00002974ffffd68c0000791a;
    assign coff[794 ] = 256'hfffff7f4ffff804100007fbffffff7f40000080c00007fbfffff80410000080c;
    assign coff[795 ] = 256'hffffab5c00006005ffff9ffbffffab5c000054a4ffff9ffb00006005000054a4;
    assign coff[796 ] = 256'h00004048ffff915000006eb000004048ffffbfb800006eb0ffff9150ffffbfb8;
    assign coff[797 ] = 256'hffff8447000020d0ffffdf30ffff844700007bb9ffffdf30000020d000007bb9;
    assign coff[798 ] = 256'hffffb257ffff9a40000065c0ffffb25700004da9000065c0ffff9a4000004da9;
    assign coff[799 ] = 256'hffffeef800007eddffff8123ffffeef800001108ffff812300007edd00001108;
    assign coff[800 ] = 256'h00007f83fffff4d300000b2d00007f83ffff807d00000b2dfffff4d3ffff807d;
    assign coff[801 ] = 256'hffff9defffffadbd00005243ffff9def0000621100005243ffffadbd00006211;
    assign coff[802 ] = 256'h00002678ffff85eb00007a1500002678ffffd98800007a15ffff85ebffffd988;
    assign coff[803 ] = 256'hffff8e7900003b20ffffc4e0ffff8e7900007187ffffc4e000003b2000007187;
    assign coff[804 ] = 256'h000063d0ffffafdd00005023000063d0ffff9c3000005023ffffafddffff9c30;
    assign coff[805 ] = 256'hffff80c2fffff21600000deaffff80c200007f3e00000deafffff21600007f3e;
    assign coff[806 ] = 256'hffffdc29ffff851f00007ae1ffffdc29000023d700007ae1ffff851f000023d7;
    assign coff[807 ] = 256'hffffc2740000703bffff8fc5ffffc27400003d8cffff8fc50000703b00003d8c;
    assign coff[808 ] = 256'h000076c7ffffd04a00002fb6000076c7ffff893900002fb6ffffd04affff8939;
    assign coff[809 ] = 256'hffff8a47ffffcdc000003240ffff8a47000075b900003240ffffcdc0000075b9;
    assign coff[810 ] = 256'h00000160ffff800200007ffe00000160fffffea000007ffeffff8002fffffea0;
    assign coff[811 ] = 256'hffffa48600005988ffffa678ffffa48600005b7affffa6780000598800005b7a;
    assign coff[812 ] = 256'h00004840ffff9657000069a900004840ffffb7c0000069a9ffff9657ffffb7c0;
    assign coff[813 ] = 256'hffff82330000179fffffe861ffff823300007dcdffffe8610000179f00007dcd;
    assign coff[814 ] = 256'hffffba09ffff94d000006b30ffffba09000045f700006b30ffff94d0000045f7;
    assign coff[815 ] = 256'hffffe5af00007d44ffff82bcffffe5af00001a51ffff82bc00007d4400001a51;
    assign coff[816 ] = 256'h00007c7effffe23c00001dc400007c7effff838200001dc4ffffe23cffff8382;
    assign coff[817 ] = 256'hffff92ecffffbd05000042fbffff92ec00006d14000042fbffffbd0500006d14;
    assign coff[818 ] = 256'h00001424ffff819800007e6800001424ffffebdc00007e68ffff8198ffffebdc;
    assign coff[819 ] = 256'hffff986000004b24ffffb4dcffff9860000067a0ffffb4dc00004b24000067a0;
    assign coff[820 ] = 256'h000056f9ffffa21600005dea000056f9ffffa90700005deaffffa216ffffa907;
    assign coff[821 ] = 256'hffff8018000004e8fffffb18ffff801800007fe8fffffb18000004e800007fe8;
    assign coff[822 ] = 256'hffffca85ffff8bb50000744bffffca850000357b0000744bffff8bb50000357b;
    assign coff[823 ] = 256'hffffd3960000780cffff87f4ffffd39600002c6affff87f40000780c00002c6a;
    assign coff[824 ] = 256'h00006e7dffffbf610000409f00006e7dffff91830000409fffffbf61ffff9183;
    assign coff[825 ] = 256'hffff842dffffdf910000206fffff842d00007bd30000206fffffdf9100007bd3;
    assign coff[826 ] = 256'hffffee94ffff813100007ecfffffee940000116c00007ecfffff81310000116c;
    assign coff[827 ] = 256'hffffb2a7000065fcffff9a04ffffb2a700004d59ffff9a04000065fc00004d59;
    assign coff[828 ] = 256'h000037f7ffff8ce20000731e000037f7ffffc8090000731effff8ce2ffffc809;
    assign coff[829 ] = 256'hffff8707000029d3ffffd62dffff8707000078f9ffffd62d000029d3000078f9;
    assign coff[830 ] = 256'hffffab10ffffa03e00005fc2ffffab10000054f000005fc2ffffa03e000054f0;
    assign coff[831 ] = 256'hfffff85900007fc5ffff803bfffff859000007a7ffff803b00007fc5000007a7;
    assign coff[832 ] = 256'h00007fd6fffff9860000067a00007fd6ffff802a0000067afffff986ffff802a;
    assign coff[833 ] = 256'hffffa107ffffaa30000055d0ffffa10700005ef9000055d0ffffaa3000005ef9;
    assign coff[834 ] = 256'h00002af0ffff876b0000789500002af0ffffd51000007895ffff876bffffd510;
    assign coff[835 ] = 256'hffff8c60000036e8ffffc918ffff8c60000073a0ffffc918000036e8000073a0;
    assign coff[836 ] = 256'h000066b2ffffb39800004c68000066b2ffff994e00004c68ffffb398ffff994e;
    assign coff[837 ] = 256'hffff815bffffed6a00001296ffff815b00007ea500001296ffffed6a00007ea5;
    assign coff[838 ] = 256'hffffe0b5ffff83e200007c1effffe0b500001f4b00007c1effff83e200001f4b;
    assign coff[839 ] = 256'hffffbe5d00006de4ffff921cffffbe5d000041a3ffff921c00006de4000041a3;
    assign coff[840 ] = 256'h00007874ffffd4b100002b4f00007874ffff878c00002b4fffffd4b1ffff878c;
    assign coff[841 ] = 256'hffff8c35ffffc9730000368dffff8c35000073cb0000368dffffc973000073cb;
    assign coff[842 ] = 256'h00000616ffff802500007fdb00000616fffff9ea00007fdbffff8025fffff9ea;
    assign coff[843 ] = 256'hffffa14a0000561bffffa9e5ffffa14a00005eb6ffffa9e50000561b00005eb6;
    assign coff[844 ] = 256'h00004c17ffff9913000066ed00004c17ffffb3e9000066edffff9913ffffb3e9;
    assign coff[845 ] = 256'hffff816a000012faffffed06ffff816a00007e96ffffed06000012fa00007e96;
    assign coff[846 ] = 256'hffffbe07ffff925000006db0ffffbe07000041f900006db0ffff9250000041f9;
    assign coff[847 ] = 256'hffffe11700007c36ffff83caffffe11700001ee9ffff83ca00007c3600001ee9;
    assign coff[848 ] = 256'h00007d81ffffe6d60000192a00007d81ffff827f0000192affffe6d6ffff827f;
    assign coff[849 ] = 256'hffff9577ffffb90d000046f3ffff957700006a89000046f3ffffb90d00006a89;
    assign coff[850 ] = 256'h000018c7ffff826c00007d94000018c7ffffe73900007d94ffff826cffffe739;
    assign coff[851 ] = 256'hffff95ae00004747ffffb8b9ffff95ae00006a52ffffb8b90000474700006a52;
    assign coff[852 ] = 256'h00005a5fffffa55a00005aa600005a5fffffa5a100005aa6ffffa55affffa5a1;
    assign coff[853 ] = 256'hffff800100000032ffffffceffff800100007fffffffffce0000003200007fff;
    assign coff[854 ] = 256'hffffced6ffff89d20000762effffced60000312a0000762effff89d20000312a;
    assign coff[855 ] = 256'hffffcf3300007655ffff89abffffcf33000030cdffff89ab00007655000030cd;
    assign coff[856 ] = 256'h000070cbffffc37d00003c83000070cbffff8f3500003c83ffffc37dffff8f35;
    assign coff[857 ] = 256'hffff8574ffffdb08000024f8ffff857400007a8c000024f8ffffdb0800007a8c;
    assign coff[858 ] = 256'hfffff342ffff80a300007f5dfffff34200000cbe00007f5dffff80a300000cbe;
    assign coff[859 ] = 256'hffffaef300006312ffff9ceeffffaef30000510dffff9cee000063120000510d;
    assign coff[860 ] = 256'h00003c2affff8f06000070fa00003c2affffc3d6000070faffff8f06ffffc3d6;
    assign coff[861 ] = 256'hffff859200002558ffffdaa8ffff859200007a6effffdaa80000255800007a6e;
    assign coff[862 ] = 256'hffffaea5ffff9d2e000062d2ffffaea50000515b000062d2ffff9d2e0000515b;
    assign coff[863 ] = 256'hfffff3a600007f67ffff8099fffff3a600000c5affff809900007f6700000c5a;
    assign coff[864 ] = 256'h00007f03fffff02300000fdd00007f03ffff80fd00000fddfffff023ffff80fd;
    assign coff[865 ] = 256'hffff9af9ffffb16800004e98ffff9af90000650700004e98ffffb16800006507;
    assign coff[866 ] = 256'h000021f3ffff849600007b6a000021f3ffffde0d00007b6affff8496ffffde0d;
    assign coff[867 ] = 256'hffff90ba00003f43ffffc0bdffff90ba00006f46ffffc0bd00003f4300006f46;
    assign coff[868 ] = 256'h000060cbffffac3f000053c1000060cbffff9f35000053c1ffffac3fffff9f35;
    assign coff[869 ] = 256'hffff8055fffff6c800000938ffff805500007fab00000938fffff6c800007fab;
    assign coff[870 ] = 256'hffffd7aaffff86860000797affffd7aa000028560000797affff868600002856;
    assign coff[871 ] = 256'hffffc6a00000726cffff8d94ffffc6a000003960ffff8d940000726c00003960;
    assign coff[872 ] = 256'h000074f0ffffcbf30000340d000074f0ffff8b100000340dffffcbf3ffff8b10;
    assign coff[873 ] = 256'hffff8882ffffd21e00002de2ffff88820000777e00002de2ffffd21e0000777e;
    assign coff[874 ] = 256'hfffffcaaffff800b00007ff5fffffcaa0000035600007ff5ffff800b00000356;
    assign coff[875 ] = 256'hffffa7e200005cd7ffffa329ffffa7e20000581effffa32900005cd70000581e;
    assign coff[876 ] = 256'h00004450ffff93c100006c3f00004450ffffbbb000006c3fffff93c1ffffbbb0;
    assign coff[877 ] = 256'hffff832700001c3dffffe3c3ffff832700007cd9ffffe3c300001c3d00007cd9;
    assign coff[878 ] = 256'hffffb623ffff97760000688affffb623000049dd0000688affff9776000049dd;
    assign coff[879 ] = 256'hffffea4f00007e26ffff81daffffea4f000015b1ffff81da00007e26000015b1;
    assign coff[880 ] = 256'h00007b50ffffddac0000225400007b50ffff84b000002254ffffddacffff84b0;
    assign coff[881 ] = 256'hffff9088ffffc11400003eecffff908800006f7800003eecffffc11400006f78;
    assign coff[882 ] = 256'h00000f79ffff80f000007f1000000f79fffff08700007f10ffff80f0fffff087;
    assign coff[883 ] = 256'hffff9b3600004ee8ffffb118ffff9b36000064caffffb11800004ee8000064ca;
    assign coff[884 ] = 256'h00005375ffff9ef30000610d00005375ffffac8b0000610dffff9ef3ffffac8b;
    assign coff[885 ] = 256'hffff805d0000099dfffff663ffff805d00007fa3fffff6630000099d00007fa3;
    assign coff[886 ] = 256'hffffc646ffff8dc10000723fffffc646000039ba0000723fffff8dc1000039ba;
    assign coff[887 ] = 256'hffffd8090000799affff8666ffffd809000027f7ffff86660000799a000027f7;
    assign coff[888 ] = 256'h00006c09ffffbb5b000044a500006c09ffff93f7000044a5ffffbb5bffff93f7;
    assign coff[889 ] = 256'hffff8311ffffe42600001bdaffff831100007cef00001bdaffffe42600007cef;
    assign coff[890 ] = 256'hffffe9ecffff81eb00007e15ffffe9ec0000161400007e15ffff81eb00001614;
    assign coff[891 ] = 256'hffffb675000068c4ffff973cffffb6750000498bffff973c000068c40000498b;
    assign coff[892 ] = 256'h000033b1ffff8ae700007519000033b1ffffcc4f00007519ffff8ae7ffffcc4f;
    assign coff[893 ] = 256'hffff88a600002e40ffffd1c0ffff88a60000775affffd1c000002e400000775a;
    assign coff[894 ] = 256'hffffa799ffffa36f00005c91ffffa7990000586700005c91ffffa36f00005867;
    assign coff[895 ] = 256'hfffffd0e00007ff7ffff8009fffffd0e000002f2ffff800900007ff7000002f2;
    assign coff[896 ] = 256'h00007feffffffbe10000041f00007fefffff80110000041ffffffbe1ffff8011;
    assign coff[897 ] = 256'hffffa29fffffa8740000578cffffa29f00005d610000578cffffa87400005d61;
    assign coff[898 ] = 256'h00002d26ffff883a000077c600002d26ffffd2da000077c6ffff883affffd2da;
    assign coff[899 ] = 256'hffff8b62000034c4ffffcb3cffff8b620000749effffcb3c000034c40000749e;
    assign coff[900 ] = 256'h00006815ffffb57f00004a8100006815ffff97eb00004a81ffffb57fffff97eb;
    assign coff[901 ] = 256'hffff81b8ffffeb16000014eaffff81b800007e48000014eaffffeb1600007e48;
    assign coff[902 ] = 256'hffffe2ffffff835400007cacffffe2ff00001d0100007cacffff835400001d01;
    assign coff[903 ] = 256'hffffbc5a00006caaffff9356ffffbc5a000043a6ffff935600006caa000043a6;
    assign coff[904 ] = 256'h0000793affffd6eb000029150000793affff86c600002915ffffd6ebffff86c6;
    assign coff[905 ] = 256'hffff8d3bffffc754000038acffff8d3b000072c5000038acffffc754000072c5;
    assign coff[906 ] = 256'h00000870ffff804700007fb900000870fffff79000007fb9ffff8047fffff790;
    assign coff[907 ] = 256'hffff9fb900005459ffffaba7ffff9fb900006047ffffaba70000545900006047;
    assign coff[908 ] = 256'h00004df9ffff9a7e0000658200004df9ffffb20700006582ffff9a7effffb207;
    assign coff[909 ] = 256'hffff8116000010a4ffffef5cffff811600007eeaffffef5c000010a400007eea;
    assign coff[910 ] = 256'hffffc00fffff911e00006ee2ffffc00f00003ff100006ee2ffff911e00003ff1;
    assign coff[911 ] = 256'hffffdecf00007b9fffff8461ffffdecf00002131ffff846100007b9f00002131;
    assign coff[912 ] = 256'h00007df2ffffe926000016da00007df2ffff820e000016daffffe926ffff820e;
    assign coff[913 ] = 256'hffff96c9ffffb71a000048e6ffff96c900006937000048e6ffffb71a00006937;
    assign coff[914 ] = 256'h00001b16ffff82e600007d1a00001b16ffffe4ea00007d1affff82e6ffffe4ea;
    assign coff[915 ] = 256'hffff94630000454fffffbab1ffff946300006b9dffffbab10000454f00006b9d;
    assign coff[916 ] = 256'h00005c06ffffa708000058f800005c06ffffa3fa000058f8ffffa708ffffa3fa;
    assign coff[917 ] = 256'hffff8005fffffdd700000229ffff800500007ffb00000229fffffdd700007ffb;
    assign coff[918 ] = 256'hffffd105ffff88ef00007711ffffd10500002efb00007711ffff88ef00002efb;
    assign coff[919 ] = 256'hffffcd070000756affff8a96ffffcd07000032f9ffff8a960000756a000032f9;
    assign coff[920 ] = 256'h000071e3ffffc59300003a6d000071e3ffff8e1d00003a6dffffc593ffff8e1d;
    assign coff[921 ] = 256'hffff8628ffffd8c800002738ffff8628000079d800002738ffffd8c8000079d8;
    assign coff[922 ] = 256'hfffff59bffff806c00007f94fffff59b00000a6500007f94ffff806c00000a65;
    assign coff[923 ] = 256'hffffad2400006190ffff9e70ffffad24000052dcffff9e7000006190000052dc;
    assign coff[924 ] = 256'h00003e3cffff902600006fda00003e3cffffc1c400006fdaffff9026ffffc1c4;
    assign coff[925 ] = 256'hffff84e700002316ffffdceaffff84e700007b19ffffdcea0000231600007b19;
    assign coff[926 ] = 256'hffffb07bffff9bb30000644dffffb07b00004f850000644dffff9bb300004f85;
    assign coff[927 ] = 256'hfffff14e00007f27ffff80d9fffff14e00000eb2ffff80d900007f2700000eb2;
    assign coff[928 ] = 256'h00007f49fffff27a00000d8600007f49ffff80b700000d86fffff27affff80b7;
    assign coff[929 ] = 256'hffff9c6fffffaf8f00005071ffff9c6f0000639100005071ffffaf8f00006391;
    assign coff[930 ] = 256'h00002437ffff853b00007ac500002437ffffdbc900007ac5ffff853bffffdbc9;
    assign coff[931 ] = 256'hffff8f9500003d34ffffc2ccffff8f950000706bffffc2cc00003d340000706b;
    assign coff[932 ] = 256'h00006252ffffae0b000051f500006252ffff9dae000051f5ffffae0bffff9dae;
    assign coff[933 ] = 256'hffff8086fffff46e00000b92ffff808600007f7a00000b92fffff46e00007f7a;
    assign coff[934 ] = 256'hffffd9e8ffff85cd00007a33ffffd9e80000261800007a33ffff85cd00002618;
    assign coff[935 ] = 256'hffffc48700007158ffff8ea8ffffc48700003b79ffff8ea80000715800003b79;
    assign coff[936 ] = 256'h000075e1ffffce1c000031e4000075e1ffff8a1f000031e4ffffce1cffff8a1f;
    assign coff[937 ] = 256'hffff895fffffcfed00003013ffff895f000076a100003013ffffcfed000076a1;
    assign coff[938 ] = 256'hffffff05ffff800100007fffffffff05000000fb00007fffffff8001000000fb;
    assign coff[939 ] = 256'hffffa63000005b34ffffa4ccffffa630000059d0ffffa4cc00005b34000059d0;
    assign coff[940 ] = 256'h0000464bffff950800006af80000464bffffb9b500006af8ffff9508ffffb9b5;
    assign coff[941 ] = 256'hffff82a8000019efffffe611ffff82a800007d58ffffe611000019ef00007d58;
    assign coff[942 ] = 256'hffffb813ffff961f000069e1ffffb813000047ed000069e1ffff961f000047ed;
    assign coff[943 ] = 256'hffffe7fe00007dbaffff8246ffffe7fe00001802ffff824600007dba00001802;
    assign coff[944 ] = 256'h00007becffffdff20000200e00007becffff84140000200effffdff2ffff8414;
    assign coff[945 ] = 256'hffff91b6ffffbf0a000040f6ffff91b600006e4a000040f6ffffbf0a00006e4a;
    assign coff[946 ] = 256'h000011cfffff813f00007ec1000011cfffffee3100007ec1ffff813fffffee31;
    assign coff[947 ] = 256'hffff99c700004d09ffffb2f7ffff99c700006639ffffb2f700004d0900006639;
    assign coff[948 ] = 256'h0000553bffffa08000005f800000553bffffaac500005f80ffffa080ffffaac5;
    assign coff[949 ] = 256'hffff803500000743fffff8bdffff803500007fcbfffff8bd0000074300007fcb;
    assign coff[950 ] = 256'hffffc863ffff8cb60000734affffc8630000379d0000734affff8cb60000379d;
    assign coff[951 ] = 256'hffffd5ce000078d8ffff8728ffffd5ce00002a32ffff8728000078d800002a32;
    assign coff[952 ] = 256'h00006d48ffffbd5b000042a500006d48ffff92b8000042a5ffffbd5bffff92b8;
    assign coff[953 ] = 256'hffff839affffe1da00001e26ffff839a00007c6600001e26ffffe1da00007c66;
    assign coff[954 ] = 256'hffffec3fffff818800007e78ffffec3f000013c100007e78ffff8188000013c1;
    assign coff[955 ] = 256'hffffb48b00006764ffff989cffffb48b00004b75ffff989c0000676400004b75;
    assign coff[956 ] = 256'h000035d7ffff8bdf00007421000035d7ffffca2900007421ffff8bdfffffca29;
    assign coff[957 ] = 256'hffff87d100002c0cffffd3f4ffff87d10000782fffffd3f400002c0c0000782f;
    assign coff[958 ] = 256'hffffa951ffffa1d200005e2effffa951000056af00005e2effffa1d2000056af;
    assign coff[959 ] = 256'hfffffab300007fe4ffff801cfffffab30000054dffff801c00007fe40000054d;
    assign coff[960 ] = 256'h00007fb2fffff72c000008d400007fb2ffff804e000008d4fffff72cffff804e;
    assign coff[961 ] = 256'hffff9f77ffffabf30000540dffff9f77000060890000540dffffabf300006089;
    assign coff[962 ] = 256'h000028b6ffff86a50000795b000028b6ffffd74a0000795bffff86a5ffffd74a;
    assign coff[963 ] = 256'hffff8d6700003906ffffc6faffff8d6700007299ffffc6fa0000390600007299;
    assign coff[964 ] = 256'h00006545ffffb1b700004e4900006545ffff9abb00004e49ffffb1b7ffff9abb;
    assign coff[965 ] = 256'hffff8109ffffefbf00001041ffff810900007ef700001041ffffefbf00007ef7;
    assign coff[966 ] = 256'hffffde6effff847b00007b85ffffde6e0000219200007b85ffff847b00002192;
    assign coff[967 ] = 256'hffffc06600006f14ffff90ecffffc06600003f9affff90ec00006f1400003f9a;
    assign coff[968 ] = 256'h000077a2ffffd27c00002d84000077a2ffff885e00002d84ffffd27cffff885e;
    assign coff[969 ] = 256'hffff8b39ffffcb9700003469ffff8b39000074c700003469ffffcb97000074c7;
    assign coff[970 ] = 256'h000003bbffff800e00007ff2000003bbfffffc4500007ff2ffff800efffffc45;
    assign coff[971 ] = 256'hffffa2e4000057d5ffffa82bffffa2e400005d1cffffa82b000057d500005d1c;
    assign coff[972 ] = 256'h00004a2fffff97b00000685000004a2fffffb5d100006850ffff97b0ffffb5d1;
    assign coff[973 ] = 256'hffff81c90000154dffffeab3ffff81c900007e37ffffeab30000154d00007e37;
    assign coff[974 ] = 256'hffffbc05ffff938b00006c75ffffbc05000043fb00006c75ffff938b000043fb;
    assign coff[975 ] = 256'hffffe36100007cc2ffff833effffe36100001c9fffff833e00007cc200001c9f;
    assign coff[976 ] = 256'h00007d05ffffe48800001b7800007d05ffff82fb00001b78ffffe488ffff82fb;
    assign coff[977 ] = 256'hffff942dffffbb06000044faffff942d00006bd3000044faffffbb0600006bd3;
    assign coff[978 ] = 256'h00001677ffff81fd00007e0300001677ffffe98900007e03ffff81fdffffe989;
    assign coff[979 ] = 256'hffff970300004939ffffb6c7ffff9703000068fdffffb6c700004939000068fd;
    assign coff[980 ] = 256'h000058b0ffffa3b400005c4c000058b0ffffa75000005c4cffffa3b4ffffa750;
    assign coff[981 ] = 256'hffff80070000028dfffffd73ffff800700007ff9fffffd730000028d00007ff9;
    assign coff[982 ] = 256'hffffccabffff8abe00007542ffffccab0000335500007542ffff8abe00003355;
    assign coff[983 ] = 256'hffffd16200007736ffff88caffffd16200002e9effff88ca0000773600002e9e;
    assign coff[984 ] = 256'h00006fa9ffffc16c00003e9400006fa9ffff905700003e94ffffc16cffff9057;
    assign coff[985 ] = 256'hffff84ccffffdd4b000022b5ffff84cc00007b34000022b5ffffdd4b00007b34;
    assign coff[986 ] = 256'hfffff0ebffff80e400007f1cfffff0eb00000f1500007f1cffff80e400000f15;
    assign coff[987 ] = 256'hffffb0c90000648bffff9b75ffffb0c900004f37ffff9b750000648b00004f37;
    assign coff[988 ] = 256'h00003a13ffff8def0000721100003a13ffffc5ed00007211ffff8defffffc5ed;
    assign coff[989 ] = 256'hffff864700002797ffffd869ffff8647000079b9ffffd86900002797000079b9;
    assign coff[990 ] = 256'hffffacd7ffff9eb20000614effffacd7000053290000614effff9eb200005329;
    assign coff[991 ] = 256'hfffff5ff00007f9cffff8064fffff5ff00000a01ffff806400007f9c00000a01;
    assign coff[992 ] = 256'h00007eb3ffffedcd0000123300007eb3ffff814d00001233ffffedcdffff814d;
    assign coff[993 ] = 256'hffff998bffffb34700004cb9ffff998b0000667500004cb9ffffb34700006675;
    assign coff[994 ] = 256'h00001facffff83fb00007c0500001facffffe05400007c05ffff83fbffffe054;
    assign coff[995 ] = 256'hffff91e90000414dffffbeb3ffff91e900006e17ffffbeb30000414d00006e17;
    assign coff[996 ] = 256'h00005f3cffffaa7a0000558600005f3cffffa0c400005586ffffaa7affffa0c4;
    assign coff[997 ] = 256'hffff802ffffff922000006deffff802f00007fd1000006defffff92200007fd1;
    assign coff[998 ] = 256'hffffd56fffff8749000078b7ffffd56f00002a91000078b7ffff874900002a91;
    assign coff[999 ] = 256'hffffc8be00007375ffff8c8bffffc8be00003742ffff8c8b0000737500003742;
    assign coff[1000] = 256'h000073f6ffffc9ce00003632000073f6ffff8c0a00003632ffffc9ceffff8c0a;
    assign coff[1001] = 256'hffff87afffffd45300002badffff87af0000785100002badffffd45300007851;
    assign coff[1002] = 256'hfffffa4fffff802000007fe0fffffa4f000005b100007fe0ffff8020000005b1;
    assign coff[1003] = 256'hffffa99b00005e72ffffa18effffa99b00005665ffffa18e00005e7200005665;
    assign coff[1004] = 256'h0000424fffff928400006d7c0000424fffffbdb100006d7cffff9284ffffbdb1;
    assign coff[1005] = 256'hffff83b200001e88ffffe178ffff83b200007c4effffe17800001e8800007c4e;
    assign coff[1006] = 256'hffffb439ffff98d700006729ffffb43900004bc700006729ffff98d700004bc7;
    assign coff[1007] = 256'hffffeca300007e87ffff8179ffffeca30000135dffff817900007e870000135d;
    assign coff[1008] = 256'h00007aa8ffffdb680000249800007aa8ffff855800002498ffffdb68ffff8558;
    assign coff[1009] = 256'hffff8f65ffffc32400003cdcffff8f650000709b00003cdcffffc3240000709b;
    assign coff[1010] = 256'h00000d22ffff80ad00007f5300000d22fffff2de00007f53ffff80adfffff2de;
    assign coff[1011] = 256'hffff9caf000050bfffffaf41ffff9caf00006351ffffaf41000050bf00006351;
    assign coff[1012] = 256'h000051a8ffff9d6e00006292000051a8ffffae5800006292ffff9d6effffae58;
    assign coff[1013] = 256'hffff808f00000bf6fffff40affff808f00007f71fffff40a00000bf600007f71;
    assign coff[1014] = 256'hffffc42effff8ed60000712affffc42e00003bd20000712affff8ed600003bd2;
    assign coff[1015] = 256'hffffda4800007a51ffff85afffffda48000025b8ffff85af00007a51000025b8;
    assign coff[1016] = 256'h00006ac1ffffb9610000469f00006ac1ffff953f0000469fffffb961ffff953f;
    assign coff[1017] = 256'hffff8293ffffe6730000198dffff829300007d6d0000198dffffe67300007d6d;
    assign coff[1018] = 256'hffffe79bffff825900007da7ffffe79b0000186500007da7ffff825900001865;
    assign coff[1019] = 256'hffffb86600006a1affff95e6ffffb8660000479affff95e600006a1a0000479a;
    assign coff[1020] = 256'h00003187ffff89f80000760800003187ffffce7900007608ffff89f8ffffce79;
    assign coff[1021] = 256'hffff898500003070ffffcf90ffff89850000767bffffcf90000030700000767b;
    assign coff[1022] = 256'hffffa5e8ffffa51300005aedffffa5e800005a1800005aedffffa51300005a18;
    assign coff[1023] = 256'hffffff6900007fffffff8001ffffff6900000097ffff800100007fff00000097;
    assign coff[1024] = 256'h00007fffffffffb50000004b00007fffffff80010000004bffffffb5ffff8001;
    assign coff[1025] = 256'hffffa548ffffa5b300005a4dffffa54800005ab800005a4dffffa5b300005ab8;
    assign coff[1026] = 256'h000030b6ffff89a20000765e000030b6ffffcf4a0000765effff89a2ffffcf4a;
    assign coff[1027] = 256'hffff89db00003141ffffcebfffff89db00007625ffffcebf0000314100007625;
    assign coff[1028] = 256'h00006a44ffffb8a40000475c00006a44ffff95bc0000475cffffb8a4ffff95bc;
    assign coff[1029] = 256'hffff8267ffffe751000018afffff826700007d99000018afffffe75100007d99;
    assign coff[1030] = 256'hffffe6bdffff828400007d7cffffe6bd0000194300007d7cffff828400001943;
    assign coff[1031] = 256'hffffb92200006a97ffff9569ffffb922000046deffff956900006a97000046de;
    assign coff[1032] = 256'h00007a67ffffda900000257000007a67ffff859900002570ffffda90ffff8599;
    assign coff[1033] = 256'hffff8efaffffc3ec00003c14ffff8efa0000710600003c14ffffc3ec00007106;
    assign coff[1034] = 256'h00000c41ffff809600007f6a00000c41fffff3bf00007f6affff8096fffff3bf;
    assign coff[1035] = 256'hffff9d3e0000516effffae92ffff9d3e000062c2ffffae920000516e000062c2;
    assign coff[1036] = 256'h000050f9ffff9cde00006322000050f9ffffaf0700006322ffff9cdeffffaf07;
    assign coff[1037] = 256'hffff80a500000cd7fffff329ffff80a500007f5bfffff32900000cd700007f5b;
    assign coff[1038] = 256'hffffc367ffff8f41000070bfffffc36700003c99000070bfffff8f4100003c99;
    assign coff[1039] = 256'hffffdb2000007a93ffff856dffffdb20000024e0ffff856d00007a93000024e0;
    assign coff[1040] = 256'h00007e92ffffeced0000131300007e92ffff816e00001313ffffecedffff816e;
    assign coff[1041] = 256'hffff9904ffffb3fd00004c03ffff9904000066fc00004c03ffffb3fd000066fc;
    assign coff[1042] = 256'h00001ed1ffff83c400007c3c00001ed1ffffe12f00007c3cffff83c4ffffe12f;
    assign coff[1043] = 256'hffff925d0000420fffffbdf1ffff925d00006da3ffffbdf10000420f00006da3;
    assign coff[1044] = 256'h00005ea5ffffa9d30000562d00005ea5ffffa15b0000562dffffa9d3ffffa15b;
    assign coff[1045] = 256'hffff8024fffffa03000005fdffff802400007fdc000005fdfffffa0300007fdc;
    assign coff[1046] = 256'hffffd49affff87950000786bffffd49a00002b660000786bffff879500002b66;
    assign coff[1047] = 256'hffffc98a000073d6ffff8c2affffc98a00003676ffff8c2a000073d600003676;
    assign coff[1048] = 256'h00007396ffffc902000036fe00007396ffff8c6a000036feffffc902ffff8c6a;
    assign coff[1049] = 256'hffff8762ffffd52800002ad8ffff87620000789e00002ad8ffffd5280000789e;
    assign coff[1050] = 256'hfffff96dffff802b00007fd5fffff96d0000069300007fd5ffff802b00000693;
    assign coff[1051] = 256'hffffaa4200005f0affffa0f6ffffaa42000055beffffa0f600005f0a000055be;
    assign coff[1052] = 256'h0000418dffff920f00006df10000418dffffbe7300006df1ffff920fffffbe73;
    assign coff[1053] = 256'hffff83e800001f63ffffe09dffff83e800007c18ffffe09d00001f6300007c18;
    assign coff[1054] = 256'hffffb384ffff995d000066a3ffffb38400004c7c000066a3ffff995d00004c7c;
    assign coff[1055] = 256'hffffed8300007ea8ffff8158ffffed830000127dffff815800007ea80000127d;
    assign coff[1056] = 256'h00007fa2fffff64a000009b600007fa2ffff805e000009b6fffff64affff805e;
    assign coff[1057] = 256'hffff9ee3ffffac9e00005362ffff9ee30000611d00005362ffffac9e0000611d;
    assign coff[1058] = 256'h000027dfffff865e000079a2000027dfffffd821000079a2ffff865effffd821;
    assign coff[1059] = 256'hffff8dcd000039d0ffffc630ffff8dcd00007233ffffc630000039d000007233;
    assign coff[1060] = 256'h000064baffffb10500004efb000064baffff9b4600004efbffffb105ffff9b46;
    assign coff[1061] = 256'hffff80edfffff0a000000f60ffff80ed00007f1300000f60fffff0a000007f13;
    assign coff[1062] = 256'hffffdd94ffff84b700007b49ffffdd940000226c00007b49ffff84b70000226c;
    assign coff[1063] = 256'hffffc12a00006f84ffff907cffffc12a00003ed6ffff907c00006f8400003ed6;
    assign coff[1064] = 256'h00007751ffffd1a900002e5700007751ffff88af00002e57ffffd1a9ffff88af;
    assign coff[1065] = 256'hffff8addffffcc660000339affff8add000075230000339affffcc6600007523;
    assign coff[1066] = 256'h000002d9ffff800800007ff8000002d9fffffd2700007ff8ffff8008fffffd27;
    assign coff[1067] = 256'hffffa38000005879ffffa787ffffa38000005c80ffffa7870000587900005c80;
    assign coff[1068] = 256'h00004976ffff972e000068d200004976ffffb68a000068d2ffff972effffb68a;
    assign coff[1069] = 256'hffff81ef0000162cffffe9d4ffff81ef00007e11ffffe9d40000162c00007e11;
    assign coff[1070] = 256'hffffbb46ffff940400006bfcffffbb46000044ba00006bfcffff9404000044ba;
    assign coff[1071] = 256'hffffe43e00007cf4ffff830cffffe43e00001bc2ffff830c00007cf400001bc2;
    assign coff[1072] = 256'h00007cd3ffffe3ab00001c5500007cd3ffff832d00001c55ffffe3abffff832d;
    assign coff[1073] = 256'hffff93b4ffffbbc50000443bffff93b400006c4c0000443bffffbbc500006c4c;
    assign coff[1074] = 256'h00001598ffff81d600007e2a00001598ffffea6800007e2affff81d6ffffea68;
    assign coff[1075] = 256'hffff9785000049f2ffffb60effff97850000687bffffb60e000049f20000687b;
    assign coff[1076] = 256'h0000580cffffa31800005ce80000580cffffa7f400005ce8ffffa318ffffa7f4;
    assign coff[1077] = 256'hffff800c00000370fffffc90ffff800c00007ff4fffffc900000037000007ff4;
    assign coff[1078] = 256'hffffcbdcffff8b1a000074e6ffffcbdc00003424000074e6ffff8b1a00003424;
    assign coff[1079] = 256'hffffd23500007787ffff8879ffffd23500002dcbffff88790000778700002dcb;
    assign coff[1080] = 256'h00006f3affffc0a700003f5900006f3affff90c600003f59ffffc0a7ffff90c6;
    assign coff[1081] = 256'hffff848fffffde25000021dbffff848f00007b71000021dbffffde2500007b71;
    assign coff[1082] = 256'hfffff00affff810000007f00fffff00a00000ff600007f00ffff810000000ff6;
    assign coff[1083] = 256'hffffb17c00006517ffff9ae9ffffb17c00004e84ffff9ae90000651700004e84;
    assign coff[1084] = 256'h00003949ffff8d890000727700003949ffffc6b700007277ffff8d89ffffc6b7;
    assign coff[1085] = 256'hffff868e0000286effffd792ffff868e00007972ffffd7920000286e00007972;
    assign coff[1086] = 256'hffffac2cffff9f45000060bbffffac2c000053d4000060bbffff9f45000053d4;
    assign coff[1087] = 256'hfffff6e100007fadffff8053fffff6e10000091fffff805300007fad0000091f;
    assign coff[1088] = 256'h00007fe7fffffaff0000050100007fe7ffff801900000501fffffaffffff8019;
    assign coff[1089] = 256'hffffa205ffffa919000056e7ffffa20500005dfb000056e7ffffa91900005dfb;
    assign coff[1090] = 256'h00002c52ffff87eb0000781500002c52ffffd3ae00007815ffff87ebffffd3ae;
    assign coff[1091] = 256'hffff8bc000003592ffffca6effff8bc000007440ffffca6e0000359200007440;
    assign coff[1092] = 256'h00006791ffffb4c800004b3800006791ffff986f00004b38ffffb4c8ffff986f;
    assign coff[1093] = 256'hffff8194ffffebf50000140bffff819400007e6c0000140bffffebf500007e6c;
    assign coff[1094] = 256'hffffe223ffff838800007c78ffffe22300001ddd00007c78ffff838800001ddd;
    assign coff[1095] = 256'hffffbd1a00006d21ffff92dfffffbd1a000042e6ffff92df00006d21000042e6;
    assign coff[1096] = 256'h000078f1ffffd615000029eb000078f1ffff870f000029ebffffd615ffff870f;
    assign coff[1097] = 256'hffff8cd7ffffc81f000037e1ffff8cd700007329000037e1ffffc81f00007329;
    assign coff[1098] = 256'h0000078effff803900007fc70000078efffff87200007fc7ffff8039fffff872;
    assign coff[1099] = 256'hffffa04e00005502ffffaafeffffa04e00005fb2ffffaafe0000550200005fb2;
    assign coff[1100] = 256'h00004d45ffff99f40000660c00004d45ffffb2bb0000660cffff99f4ffffb2bb;
    assign coff[1101] = 256'hffff813400001185ffffee7bffff813400007eccffffee7b0000118500007ecc;
    assign coff[1102] = 256'hffffbf4bffff918f00006e71ffffbf4b000040b500006e71ffff918f000040b5;
    assign coff[1103] = 256'hffffdfa900007bd9ffff8427ffffdfa900002057ffff842700007bd900002057;
    assign coff[1104] = 256'h00007dc9ffffe848000017b800007dc9ffff8237000017b8ffffe848ffff8237;
    assign coff[1105] = 256'hffff9649ffffb7d40000482cffff9649000069b70000482cffffb7d4000069b7;
    assign coff[1106] = 256'h00001a39ffff82b700007d4900001a39ffffe5c700007d49ffff82b7ffffe5c7;
    assign coff[1107] = 256'hffff94de0000460cffffb9f4ffff94de00006b22ffffb9f40000460c00006b22;
    assign coff[1108] = 256'h00005b68ffffa6660000599a00005b68ffffa4980000599affffa666ffffa498;
    assign coff[1109] = 256'hffff8002fffffeb900000147ffff800200007ffe00000147fffffeb900007ffe;
    assign coff[1110] = 256'hffffd033ffff8943000076bdffffd03300002fcd000076bdffff894300002fcd;
    assign coff[1111] = 256'hffffcdd7000075c3ffff8a3dffffcdd700003229ffff8a3d000075c300003229;
    assign coff[1112] = 256'h0000717bffffc4ca00003b360000717bffff8e8500003b36ffffc4caffff8e85;
    assign coff[1113] = 256'hffff85e3ffffd9a000002660ffff85e300007a1d00002660ffffd9a000007a1d;
    assign coff[1114] = 256'hfffff4b9ffff807f00007f81fffff4b900000b4700007f81ffff807f00000b47;
    assign coff[1115] = 256'hffffadd100006221ffff9ddfffffadd10000522fffff9ddf000062210000522f;
    assign coff[1116] = 256'h00003d76ffff8fb90000704700003d76ffffc28a00007047ffff8fb9ffffc28a;
    assign coff[1117] = 256'hffff8526000023efffffdc11ffff852600007adaffffdc11000023ef00007ada;
    assign coff[1118] = 256'hffffafcaffff9c40000063c0ffffafca00005036000063c0ffff9c4000005036;
    assign coff[1119] = 256'hfffff22f00007f41ffff80bffffff22f00000dd1ffff80bf00007f4100000dd1;
    assign coff[1120] = 256'h00007f30fffff19900000e6700007f30ffff80d000000e67fffff199ffff80d0;
    assign coff[1121] = 256'hffff9be2ffffb04000004fc0ffff9be20000641e00004fc0ffffb0400000641e;
    assign coff[1122] = 256'h0000235effff84fc00007b040000235effffdca200007b04ffff84fcffffdca2;
    assign coff[1123] = 256'hffff900100003dfaffffc206ffff900100006fffffffc20600003dfa00006fff;
    assign coff[1124] = 256'h000061c0ffffad5d000052a3000061c0ffff9e40000052a3ffffad5dffff9e40;
    assign coff[1125] = 256'hffff8072fffff55000000ab0ffff807200007f8e00000ab0fffff55000007f8e;
    assign coff[1126] = 256'hffffd910ffff8611000079efffffd910000026f0000079efffff8611000026f0;
    assign coff[1127] = 256'hffffc550000071c1ffff8e3fffffc55000003ab0ffff8e3f000071c100003ab0;
    assign coff[1128] = 256'h00007588ffffcd4c000032b400007588ffff8a78000032b4ffffcd4cffff8a78;
    assign coff[1129] = 256'hffff890bffffd0bf00002f41ffff890b000076f500002f41ffffd0bf000076f5;
    assign coff[1130] = 256'hfffffe22ffff800300007ffdfffffe22000001de00007ffdffff8003000001de;
    assign coff[1131] = 256'hffffa6d200005bd2ffffa42effffa6d20000592effffa42e00005bd20000592e;
    assign coff[1132] = 256'h0000458effff948c00006b740000458effffba7200006b74ffff948cffffba72;
    assign coff[1133] = 256'hffff82d600001accffffe534ffff82d600007d2affffe53400001acc00007d2a;
    assign coff[1134] = 256'hffffb758ffff969f00006961ffffb758000048a800006961ffff969f000048a8;
    assign coff[1135] = 256'hffffe8dc00007de4ffff821cffffe8dc00001724ffff821c00007de400001724;
    assign coff[1136] = 256'h00007bb3ffffdf18000020e800007bb3ffff844d000020e8ffffdf18ffff844d;
    assign coff[1137] = 256'hffff9143ffffbfcd00004033ffff914300006ebd00004033ffffbfcd00006ebd;
    assign coff[1138] = 256'h000010efffff812000007ee0000010efffffef1100007ee0ffff8120ffffef11;
    assign coff[1139] = 256'hffff9a5000004dbdffffb243ffff9a50000065b0ffffb24300004dbd000065b0;
    assign coff[1140] = 256'h00005491ffff9fea0000601600005491ffffab6f00006016ffff9feaffffab6f;
    assign coff[1141] = 256'hffff804200000825fffff7dbffff804200007fbefffff7db0000082500007fbe;
    assign coff[1142] = 256'hffffc798ffff8d19000072e7ffffc79800003868000072e7ffff8d1900003868;
    assign coff[1143] = 256'hffffd6a400007922ffff86deffffd6a40000295cffff86de000079220000295c;
    assign coff[1144] = 256'h00006cd2ffffbc9a0000436600006cd2ffff932e00004366ffffbc9affff932e;
    assign coff[1145] = 256'hffff8365ffffe2b600001d4affff836500007c9b00001d4affffe2b600007c9b;
    assign coff[1146] = 256'hffffeb60ffff81ac00007e54ffffeb60000014a000007e54ffff81ac000014a0;
    assign coff[1147] = 256'hffffb542000067e9ffff9817ffffb54200004abeffff9817000067e900004abe;
    assign coff[1148] = 256'h00003509ffff8b810000747f00003509ffffcaf70000747fffff8b81ffffcaf7;
    assign coff[1149] = 256'hffff882000002ce0ffffd320ffff8820000077e0ffffd32000002ce0000077e0;
    assign coff[1150] = 256'hffffa8abffffa26c00005d94ffffa8ab0000575500005d94ffffa26c00005755;
    assign coff[1151] = 256'hfffffb9500007fecffff8014fffffb950000046bffff801400007fec0000046b;
    assign coff[1152] = 256'h00007ff9fffffd59000002a700007ff9ffff8007000002a7fffffd59ffff8007;
    assign coff[1153] = 256'hffffa3a3ffffa7620000589effffa3a300005c5d0000589effffa76200005c5d;
    assign coff[1154] = 256'h00002e86ffff88c10000773f00002e86ffffd17a0000773fffff88c1ffffd17a;
    assign coff[1155] = 256'hffff8ac80000336cffffcc94ffff8ac800007538ffffcc940000336c00007538;
    assign coff[1156] = 256'h000068efffffb6b30000494d000068efffff97110000494dffffb6b3ffff9711;
    assign coff[1157] = 256'hffff81f8ffffe9a20000165effff81f800007e080000165effffe9a200007e08;
    assign coff[1158] = 256'hffffe46fffff830100007cffffffe46f00001b9100007cffffff830100001b91;
    assign coff[1159] = 256'hffffbb1b00006be1ffff941fffffbb1b000044e5ffff941f00006be1000044e5;
    assign coff[1160] = 256'h000079b1ffffd851000027af000079b1ffff864f000027afffffd851ffff864f;
    assign coff[1161] = 256'hffff8de4ffffc603000039fdffff8de40000721c000039fdffffc6030000721c;
    assign coff[1162] = 256'h000009e8ffff806200007f9e000009e8fffff61800007f9effff8062fffff618;
    assign coff[1163] = 256'hffff9ec20000533cffffacc4ffff9ec20000613effffacc40000533c0000613e;
    assign coff[1164] = 256'h00004f23ffff9b650000649b00004f23ffffb0dd0000649bffff9b65ffffb0dd;
    assign coff[1165] = 256'hffff80e700000f2efffff0d2ffff80e700007f19fffff0d200000f2e00007f19;
    assign coff[1166] = 256'hffffc156ffff906300006f9dffffc15600003eaa00006f9dffff906300003eaa;
    assign coff[1167] = 256'hffffdd6300007b3bffff84c5ffffdd630000229dffff84c500007b3b0000229d;
    assign coff[1168] = 256'h00007e33ffffea9a0000156600007e33ffff81cd00001566ffffea9affff81cd;
    assign coff[1169] = 256'hffff97a2ffffb5e500004a1bffff97a20000685e00004a1bffffb5e50000685e;
    assign coff[1170] = 256'h00001c86ffff833800007cc800001c86ffffe37a00007cc8ffff8338ffffe37a;
    assign coff[1171] = 256'hffff939900004411ffffbbefffff939900006c67ffffbbef0000441100006c67;
    assign coff[1172] = 256'h00005d0bffffa818000057e800005d0bffffa2f5000057e8ffffa818ffffa2f5;
    assign coff[1173] = 256'hffff800dfffffc5e000003a2ffff800d00007ff3000003a2fffffc5e00007ff3;
    assign coff[1174] = 256'hffffd264ffff886700007799ffffd26400002d9c00007799ffff886700002d9c;
    assign coff[1175] = 256'hffffcbae000074d2ffff8b2effffcbae00003452ffff8b2e000074d200003452;
    assign coff[1176] = 256'h0000728dffffc6e30000391d0000728dffff8d730000391dffffc6e3ffff8d73;
    assign coff[1177] = 256'hffff869effffd7620000289effff869e000079620000289effffd76200007962;
    assign coff[1178] = 256'hfffff713ffff805000007fb0fffff713000008ed00007fb0ffff8050000008ed;
    assign coff[1179] = 256'hffffac060000609affff9f66ffffac06000053faffff9f660000609a000053fa;
    assign coff[1180] = 256'h00003f85ffff90df00006f2100003f85ffffc07b00006f21ffff90dfffffc07b;
    assign coff[1181] = 256'hffff8482000021aaffffde56ffff848200007b7effffde56000021aa00007b7e;
    assign coff[1182] = 256'hffffb1a3ffff9aca00006536ffffb1a300004e5d00006536ffff9aca00004e5d;
    assign coff[1183] = 256'hffffefd800007efaffff8106ffffefd800001028ffff810600007efa00001028;
    assign coff[1184] = 256'h00007f6efffff3f100000c0f00007f6effff809200000c0ffffff3f1ffff8092;
    assign coff[1185] = 256'hffff9d5effffae6b00005195ffff9d5e000062a200005195ffffae6b000062a2;
    assign coff[1186] = 256'h000025a0ffff85a800007a58000025a0ffffda6000007a58ffff85a8ffffda60;
    assign coff[1187] = 256'hffff8ee200003be8ffffc418ffff8ee20000711effffc41800003be80000711e;
    assign coff[1188] = 256'h00006342ffffaf2d000050d300006342ffff9cbe000050d3ffffaf2dffff9cbe;
    assign coff[1189] = 256'hffff80aafffff2f700000d09ffff80aa00007f5600000d09fffff2f700007f56;
    assign coff[1190] = 256'hffffdb50ffff855f00007aa1ffffdb50000024b000007aa1ffff855f000024b0;
    assign coff[1191] = 256'hffffc33b000070a7ffff8f59ffffc33b00003cc5ffff8f59000070a700003cc5;
    assign coff[1192] = 256'h00007672ffffcf780000308800007672ffff898e00003088ffffcf78ffff898e;
    assign coff[1193] = 256'hffff89efffffce9000003170ffff89ef0000761100003170ffffce9000007611;
    assign coff[1194] = 256'h0000007effff800100007fff0000007effffff8200007fffffff8001ffffff82;
    assign coff[1195] = 256'hffffa52500005a29ffffa5d7ffffa52500005adbffffa5d700005a2900005adb;
    assign coff[1196] = 256'h00004785ffff95d800006a2800004785ffffb87b00006a28ffff95d8ffffb87b;
    assign coff[1197] = 256'hffff825d0000187dffffe783ffff825d00007da3ffffe7830000187d00007da3;
    assign coff[1198] = 256'hffffb94cffff954d00006ab3ffffb94c000046b400006ab3ffff954d000046b4;
    assign coff[1199] = 256'hffffe68c00007d72ffff828effffe68c00001974ffff828e00007d7200001974;
    assign coff[1200] = 256'h00007c48ffffe16000001ea000007c48ffff83b800001ea0ffffe160ffff83b8;
    assign coff[1201] = 256'hffff9277ffffbdc60000423affff927700006d890000423affffbdc600006d89;
    assign coff[1202] = 256'h00001344ffff817500007e8b00001344ffffecbc00007e8bffff8175ffffecbc;
    assign coff[1203] = 256'hffff98e600004bdbffffb425ffff98e60000671affffb42500004bdb0000671a;
    assign coff[1204] = 256'h00005653ffffa17d00005e8300005653ffffa9ad00005e83ffffa17dffffa9ad;
    assign coff[1205] = 256'hffff8022000005cafffffa36ffff802200007fdefffffa36000005ca00007fde;
    assign coff[1206] = 256'hffffc9b8ffff8c15000073ebffffc9b800003648000073ebffff8c1500003648;
    assign coff[1207] = 256'hffffd46b0000785affff87a6ffffd46b00002b95ffff87a60000785a00002b95;
    assign coff[1208] = 256'h00006e0affffbe9e0000416200006e0affff91f600004162ffffbe9effff91f6;
    assign coff[1209] = 256'hffff83f5ffffe06c00001f94ffff83f500007c0b00001f94ffffe06c00007c0b;
    assign coff[1210] = 256'hffffedb4ffff815000007eb0ffffedb40000124c00007eb0ffff81500000124c;
    assign coff[1211] = 256'hffffb35b00006684ffff997cffffb35b00004ca5ffff997c0000668400004ca5;
    assign coff[1212] = 256'h0000372cffff8c80000073800000372cffffc8d400007380ffff8c80ffffc8d4;
    assign coff[1213] = 256'hffff875100002aa9ffffd557ffff8751000078afffffd55700002aa9000078af;
    assign coff[1214] = 256'hffffaa68ffffa0d400005f2cffffaa680000559800005f2cffffa0d400005598;
    assign coff[1215] = 256'hfffff93b00007fd2ffff802efffff93b000006c5ffff802e00007fd2000006c5;
    assign coff[1216] = 256'h00007fcafffff8a40000075c00007fcaffff80360000075cfffff8a4ffff8036;
    assign coff[1217] = 256'hffffa070ffffaad800005528ffffa07000005f9000005528ffffaad800005f90;
    assign coff[1218] = 256'h00002a1bffff871f000078e100002a1bffffd5e5000078e1ffff871fffffd5e5;
    assign coff[1219] = 256'hffff8cc1000037b4ffffc84cffff8cc10000733fffffc84c000037b40000733f;
    assign coff[1220] = 256'h0000662affffb2e300004d1d0000662affff99d600004d1dffffb2e3ffff99d6;
    assign coff[1221] = 256'hffff813bffffee4a000011b6ffff813b00007ec5000011b6ffffee4a00007ec5;
    assign coff[1222] = 256'hffffdfdaffff841a00007be6ffffdfda0000202600007be6ffff841a00002026;
    assign coff[1223] = 256'hffffbf2000006e57ffff91a9ffffbf20000040e0ffff91a900006e57000040e0;
    assign coff[1224] = 256'h00007826ffffd3dd00002c2300007826ffff87da00002c23ffffd3ddffff87da;
    assign coff[1225] = 256'hffff8bd5ffffca40000035c0ffff8bd50000742b000035c0ffffca400000742b;
    assign coff[1226] = 256'h00000534ffff801b00007fe500000534fffffacc00007fe5ffff801bfffffacc;
    assign coff[1227] = 256'hffffa1e3000056c2ffffa93effffa1e300005e1dffffa93e000056c200005e1d;
    assign coff[1228] = 256'h00004b61ffff988d0000677300004b61ffffb49f00006773ffff988dffffb49f;
    assign coff[1229] = 256'hffff818c000013d9ffffec27ffff818c00007e74ffffec27000013d900007e74;
    assign coff[1230] = 256'hffffbd45ffff92c500006d3bffffbd45000042bb00006d3bffff92c5000042bb;
    assign coff[1231] = 256'hffffe1f200007c6cffff8394ffffe1f200001e0effff839400007c6c00001e0e;
    assign coff[1232] = 256'h00007d53ffffe5f800001a0800007d53ffff82ad00001a08ffffe5f8ffff82ad;
    assign coff[1233] = 256'hffff94faffffb9ca00004636ffff94fa00006b0600004636ffffb9ca00006b06;
    assign coff[1234] = 256'h000017e9ffff824100007dbf000017e9ffffe81700007dbfffff8241ffffe817;
    assign coff[1235] = 256'hffff962d00004802ffffb7feffff962d000069d3ffffb7fe00004802000069d3;
    assign coff[1236] = 256'h000059beffffa4bb00005b45000059beffffa64200005b45ffffa4bbffffa642;
    assign coff[1237] = 256'hffff800100000114fffffeecffff800100007ffffffffeec0000011400007fff;
    assign coff[1238] = 256'hffffce05ffff8a29000075d7ffffce05000031fb000075d7ffff8a29000031fb;
    assign coff[1239] = 256'hffffd004000076aaffff8956ffffd00400002ffcffff8956000076aa00002ffc;
    assign coff[1240] = 256'h0000705fffffc2b600003d4a0000705fffff8fa100003d4affffc2b6ffff8fa1;
    assign coff[1241] = 256'hffff8534ffffdbe10000241fffff853400007acc0000241fffffdbe100007acc;
    assign coff[1242] = 256'hfffff261ffff80ba00007f46fffff26100000d9f00007f46ffff80ba00000d9f;
    assign coff[1243] = 256'hffffafa3000063a0ffff9c60ffffafa30000505dffff9c60000063a00000505d;
    assign coff[1244] = 256'h00003b62ffff8e9c0000716400003b62ffffc49e00007164ffff8e9cffffc49e;
    assign coff[1245] = 256'hffff85d400002630ffffd9d0ffff85d400007a2cffffd9d00000263000007a2c;
    assign coff[1246] = 256'hffffadf7ffff9dbe00006242ffffadf70000520900006242ffff9dbe00005209;
    assign coff[1247] = 256'hfffff48700007f7cffff8084fffff48700000b79ffff808400007f7c00000b79;
    assign coff[1248] = 256'h00007ee7ffffef43000010bd00007ee7ffff8119000010bdffffef43ffff8119;
    assign coff[1249] = 256'hffff9a6effffb21b00004de5ffff9a6e0000659200004de5ffffb21b00006592;
    assign coff[1250] = 256'h00002119ffff845a00007ba600002119ffffdee700007ba6ffff845affffdee7;
    assign coff[1251] = 256'hffff912a00004007ffffbff9ffff912a00006ed6ffffbff90000400700006ed6;
    assign coff[1252] = 256'h00006037ffffab940000546c00006037ffff9fc90000546cffffab94ffff9fc9;
    assign coff[1253] = 256'hffff8046fffff7a900000857ffff804600007fba00000857fffff7a900007fba;
    assign coff[1254] = 256'hffffd6d3ffff86ce00007932ffffd6d30000292d00007932ffff86ce0000292d;
    assign coff[1255] = 256'hffffc76b000072d0ffff8d30ffffc76b00003895ffff8d30000072d000003895;
    assign coff[1256] = 256'h00007494ffffcb25000034db00007494ffff8b6c000034dbffffcb25ffff8b6c;
    assign coff[1257] = 256'hffff8831ffffd2f100002d0fffff8831000077cf00002d0fffffd2f1000077cf;
    assign coff[1258] = 256'hfffffbc7ffff801200007feefffffbc70000043900007feeffff801200000439;
    assign coff[1259] = 256'hffffa88600005d72ffffa28effffa8860000577affffa28e00005d720000577a;
    assign coff[1260] = 256'h00004391ffff934900006cb700004391ffffbc6f00006cb7ffff9349ffffbc6f;
    assign coff[1261] = 256'hffff835a00001d19ffffe2e7ffff835a00007ca6ffffe2e700001d1900007ca6;
    assign coff[1262] = 256'hffffb56bffff97fa00006806ffffb56b00004a9500006806ffff97fa00004a95;
    assign coff[1263] = 256'hffffeb2f00007e4cffff81b4ffffeb2f000014d1ffff81b400007e4c000014d1;
    assign coff[1264] = 256'h00007b12ffffdcd20000232e00007b12ffff84ee0000232effffdcd2ffff84ee;
    assign coff[1265] = 256'hffff901affffc1da00003e26ffff901a00006fe600003e26ffffc1da00006fe6;
    assign coff[1266] = 256'h00000e99ffff80d600007f2a00000e99fffff16700007f2affff80d6fffff167;
    assign coff[1267] = 256'hffff9bc200004f99ffffb067ffff9bc20000643effffb06700004f990000643e;
    assign coff[1268] = 256'h000052c9ffff9e60000061a0000052c9ffffad37000061a0ffff9e60ffffad37;
    assign coff[1269] = 256'hffff806e00000a7efffff582ffff806e00007f92fffff58200000a7e00007f92;
    assign coff[1270] = 256'hffffc57dffff8e28000071d8ffffc57d00003a83000071d8ffff8e2800003a83;
    assign coff[1271] = 256'hffffd8e0000079e0ffff8620ffffd8e000002720ffff8620000079e000002720;
    assign coff[1272] = 256'h00006b8fffffba9c0000456400006b8fffff947100004564ffffba9cffff9471;
    assign coff[1273] = 256'hffff82e1ffffe50200001afeffff82e100007d1f00001afeffffe50200007d1f;
    assign coff[1274] = 256'hffffe90effff821300007dedffffe90e000016f200007dedffff8213000016f2;
    assign coff[1275] = 256'hffffb72f00006945ffff96bbffffb72f000048d1ffff96bb00006945000048d1;
    assign coff[1276] = 256'h000032e2ffff8a8c00007574000032e2ffffcd1e00007574ffff8a8cffffcd1e;
    assign coff[1277] = 256'hffff88f800002f13ffffd0edffff88f800007708ffffd0ed00002f1300007708;
    assign coff[1278] = 256'hffffa6f6ffffa40b00005bf5ffffa6f60000590a00005bf5ffffa40b0000590a;
    assign coff[1279] = 256'hfffffdf000007ffcffff8004fffffdf000000210ffff800400007ffc00000210;
    assign coff[1280] = 256'h00007ffefffffe870000017900007ffeffff800200000179fffffe87ffff8002;
    assign coff[1281] = 256'hffffa474ffffa68a00005976ffffa47400005b8c00005976ffffa68a00005b8c;
    assign coff[1282] = 256'h00002f9fffff8930000076d000002f9fffffd061000076d0ffff8930ffffd061;
    assign coff[1283] = 256'hffff8a5100003257ffffcda9ffff8a51000075afffffcda900003257000075af;
    assign coff[1284] = 256'h0000699affffb7ab000048550000699affff966600004855ffffb7abffff9666;
    assign coff[1285] = 256'hffff822effffe87900001787ffff822e00007dd200001787ffffe87900007dd2;
    assign coff[1286] = 256'hffffe596ffff82c100007d3fffffe59600001a6a00007d3fffff82c100001a6a;
    assign coff[1287] = 256'hffffba1e00006b3dffff94c3ffffba1e000045e2ffff94c300006b3d000045e2;
    assign coff[1288] = 256'h00007a0effffd9700000269000007a0effff85f200002690ffffd970ffff85f2;
    assign coff[1289] = 256'hffff8e6dffffc4f700003b09ffff8e6d0000719300003b09ffffc4f700007193;
    assign coff[1290] = 256'h00000b14ffff807b00007f8500000b14fffff4ec00007f85ffff807bfffff4ec;
    assign coff[1291] = 256'hffff9dff00005256ffffadaaffff9dff00006201ffffadaa0000525600006201;
    assign coff[1292] = 256'h0000500fffff9c21000063df0000500fffffaff1000063dfffff9c21ffffaff1;
    assign coff[1293] = 256'hffff80c500000e03fffff1fdffff80c500007f3bfffff1fd00000e0300007f3b;
    assign coff[1294] = 256'hffffc25effff8fd10000702fffffc25e00003da20000702fffff8fd100003da2;
    assign coff[1295] = 256'hffffdc4100007ae8ffff8518ffffdc41000023bfffff851800007ae8000023bf;
    assign coff[1296] = 256'h00007e64ffffebc30000143d00007e64ffff819c0000143dffffebc3ffff819c;
    assign coff[1297] = 256'hffff9852ffffb4f000004b10ffff9852000067ae00004b10ffffb4f0000067ae;
    assign coff[1298] = 256'h00001dacffff837d00007c8300001dacffffe25400007c83ffff837dffffe254;
    assign coff[1299] = 256'hffff92fa00004310ffffbcf0ffff92fa00006d06ffffbcf00000431000006d06;
    assign coff[1300] = 256'h00005dd9ffffa8f40000570c00005dd9ffffa2270000570cffffa8f4ffffa227;
    assign coff[1301] = 256'hffff8017fffffb31000004cfffff801700007fe9000004cffffffb3100007fe9;
    assign coff[1302] = 256'hffffd37fffff87fd00007803ffffd37f00002c8100007803ffff87fd00002c81;
    assign coff[1303] = 256'hffffca9c00007455ffff8babffffca9c00003564ffff8bab0000745500003564;
    assign coff[1304] = 256'h00007313ffffc7f20000380e00007313ffff8ced0000380effffc7f2ffff8ced;
    assign coff[1305] = 256'hffff86ffffffd644000029bcffff86ff00007901000029bcffffd64400007901;
    assign coff[1306] = 256'hfffff840ffff803c00007fc4fffff840000007c000007fc4ffff803c000007c0;
    assign coff[1307] = 256'hffffab2300005fd3ffffa02dffffab23000054ddffffa02d00005fd3000054dd;
    assign coff[1308] = 256'h0000408affff917600006e8a0000408affffbf7600006e8affff9176ffffbf76;
    assign coff[1309] = 256'hffff843400002087ffffdf79ffff843400007bccffffdf790000208700007bcc;
    assign coff[1310] = 256'hffffb293ffff9a13000065edffffb29300004d6d000065edffff9a1300004d6d;
    assign coff[1311] = 256'hffffeead00007ed3ffff812dffffeead00001153ffff812d00007ed300001153;
    assign coff[1312] = 256'h00007f89fffff51e00000ae200007f89ffff807700000ae2fffff51effff8077;
    assign coff[1313] = 256'hffff9e1fffffad840000527cffff9e1f000061e10000527cffffad84000061e1;
    assign coff[1314] = 256'h000026c0ffff8602000079fe000026c0ffffd940000079feffff8602ffffd940;
    assign coff[1315] = 256'hffff8e5600003addffffc523ffff8e56000071aaffffc52300003add000071aa;
    assign coff[1316] = 256'h000063ffffffb01800004fe8000063ffffff9c0100004fe8ffffb018ffff9c01;
    assign coff[1317] = 256'hffff80cafffff1cb00000e35ffff80ca00007f3600000e35fffff1cb00007f36;
    assign coff[1318] = 256'hffffdc72ffff850a00007af6ffffdc720000238e00007af6ffff850a0000238e;
    assign coff[1319] = 256'hffffc23200007017ffff8fe9ffffc23200003dceffff8fe90000701700003dce;
    assign coff[1320] = 256'h000076e3ffffd09000002f70000076e3ffff891d00002f70ffffd090ffff891d;
    assign coff[1321] = 256'hffff8a64ffffcd7b00003285ffff8a640000759c00003285ffffcd7b0000759c;
    assign coff[1322] = 256'h000001abffff800300007ffd000001abfffffe5500007ffdffff8003fffffe55;
    assign coff[1323] = 256'hffffa45100005952ffffa6aeffffa45100005bafffffa6ae0000595200005baf;
    assign coff[1324] = 256'h0000487fffff96820000697e0000487fffffb7810000697effff9682ffffb781;
    assign coff[1325] = 256'hffff822500001755ffffe8abffff822500007ddbffffe8ab0000175500007ddb;
    assign coff[1326] = 256'hffffba48ffff94a700006b59ffffba48000045b800006b59ffff94a7000045b8;
    assign coff[1327] = 256'hffffe56500007d34ffff82ccffffe56500001a9bffff82cc00007d3400001a9b;
    assign coff[1328] = 256'h00007c8fffffe28500001d7b00007c8fffff837100001d7bffffe285ffff8371;
    assign coff[1329] = 256'hffff9314ffffbcc50000433bffff931400006cec0000433bffffbcc500006cec;
    assign coff[1330] = 256'h0000146effff81a400007e5c0000146effffeb9200007e5cffff81a4ffffeb92;
    assign coff[1331] = 256'hffff983400004ae7ffffb519ffff9834000067ccffffb51900004ae7000067cc;
    assign coff[1332] = 256'h00005730ffffa24900005db700005730ffffa8d000005db7ffffa249ffffa8d0;
    assign coff[1333] = 256'hffff80150000049dfffffb63ffff801500007febfffffb630000049d00007feb;
    assign coff[1334] = 256'hffffcac9ffff8b960000746affffcac9000035370000746affff8b9600003537;
    assign coff[1335] = 256'hffffd34f000077f2ffff880effffd34f00002cb1ffff880e000077f200002cb1;
    assign coff[1336] = 256'h00006ea3ffffbfa20000405e00006ea3ffff915d0000405effffbfa2ffff915d;
    assign coff[1337] = 256'hffff8441ffffdf48000020b8ffff844100007bbf000020b8ffffdf4800007bbf;
    assign coff[1338] = 256'hffffeedfffff812700007ed9ffffeedf0000112100007ed9ffff812700001121;
    assign coff[1339] = 256'hffffb26b000065cfffff9a31ffffb26b00004d95ffff9a31000065cf00004d95;
    assign coff[1340] = 256'h0000383bffff8d03000072fd0000383bffffc7c5000072fdffff8d03ffffc7c5;
    assign coff[1341] = 256'hffff86ee0000298cffffd674ffff86ee00007912ffffd6740000298c00007912;
    assign coff[1342] = 256'hffffab49ffffa00c00005ff4ffffab49000054b700005ff4ffffa00c000054b7;
    assign coff[1343] = 256'hfffff80e00007fc1ffff803ffffff80e000007f2ffff803f00007fc1000007f2;
    assign coff[1344] = 256'h00007fdafffff9d10000062f00007fdaffff80260000062ffffff9d1ffff8026;
    assign coff[1345] = 256'hffffa139ffffa9f800005608ffffa13900005ec700005608ffffa9f800005ec7;
    assign coff[1346] = 256'h00002b37ffff87840000787c00002b37ffffd4c90000787cffff8784ffffd4c9;
    assign coff[1347] = 256'hffff8c3f000036a3ffffc95dffff8c3f000073c1ffffc95d000036a3000073c1;
    assign coff[1348] = 256'h000066deffffb3d400004c2c000066deffff992200004c2cffffb3d4ffff9922;
    assign coff[1349] = 256'hffff8166ffffed1f000012e1ffff816600007e9a000012e1ffffed1f00007e9a;
    assign coff[1350] = 256'hffffe0feffff83d000007c30ffffe0fe00001f0200007c30ffff83d000001f02;
    assign coff[1351] = 256'hffffbe1c00006dbdffff9243ffffbe1c000041e4ffff924300006dbd000041e4;
    assign coff[1352] = 256'h0000788dffffd4f800002b080000788dffff877300002b08ffffd4f8ffff8773;
    assign coff[1353] = 256'hffff8c55ffffc92f000036d1ffff8c55000073ab000036d1ffffc92f000073ab;
    assign coff[1354] = 256'h00000661ffff802900007fd700000661fffff99f00007fd7ffff8029fffff99f;
    assign coff[1355] = 256'hffffa118000055e3ffffaa1dffffa11800005ee8ffffaa1d000055e300005ee8;
    assign coff[1356] = 256'h00004c54ffff993f000066c100004c54ffffb3ac000066c1ffff993fffffb3ac;
    assign coff[1357] = 256'hffff815f000012afffffed51ffff815f00007ea1ffffed51000012af00007ea1;
    assign coff[1358] = 256'hffffbe47ffff922900006dd7ffffbe47000041b900006dd7ffff9229000041b9;
    assign coff[1359] = 256'hffffe0ce00007c24ffff83dcffffe0ce00001f32ffff83dc00007c2400001f32;
    assign coff[1360] = 256'h00007d8fffffe720000018e000007d8fffff8271000018e0ffffe720ffff8271;
    assign coff[1361] = 256'hffff95a0ffffb8ce00004732ffff95a000006a6000004732ffffb8ce00006a60;
    assign coff[1362] = 256'h00001911ffff827b00007d8500001911ffffe6ef00007d85ffff827bffffe6ef;
    assign coff[1363] = 256'hffff958400004708ffffb8f8ffff958400006a7cffffb8f80000470800006a7c;
    assign coff[1364] = 256'h00005a94ffffa58f00005a7100005a94ffffa56c00005a71ffffa58fffffa56c;
    assign coff[1365] = 256'hffff8001ffffffe700000019ffff800100007fff00000019ffffffe700007fff;
    assign coff[1366] = 256'hffffcf1bffff89b50000764bffffcf1b000030e50000764bffff89b5000030e5;
    assign coff[1367] = 256'hffffceed00007638ffff89c8ffffceed00003113ffff89c80000763800003113;
    assign coff[1368] = 256'h000070efffffc3bf00003c41000070efffff8f1100003c41ffffc3bfffff8f11;
    assign coff[1369] = 256'hffff858affffdac000002540ffff858a00007a7600002540ffffdac000007a76;
    assign coff[1370] = 256'hfffff38dffff809b00007f65fffff38d00000c7300007f65ffff809b00000c73;
    assign coff[1371] = 256'hffffaeb9000062e2ffff9d1effffaeb900005147ffff9d1e000062e200005147;
    assign coff[1372] = 256'h00003c6dffff8f29000070d700003c6dffffc393000070d7ffff8f29ffffc393;
    assign coff[1373] = 256'hffff857c00002510ffffdaf0ffff857c00007a84ffffdaf00000251000007a84;
    assign coff[1374] = 256'hffffaee0ffff9cfe00006302ffffaee00000512000006302ffff9cfe00005120;
    assign coff[1375] = 256'hfffff35b00007f60ffff80a0fffff35b00000ca5ffff80a000007f6000000ca5;
    assign coff[1376] = 256'h00007f0dfffff06e00000f9200007f0dffff80f300000f92fffff06effff80f3;
    assign coff[1377] = 256'hffff9b27ffffb12c00004ed4ffff9b27000064d900004ed4ffffb12c000064d9;
    assign coff[1378] = 256'h0000223cffff84aa00007b560000223cffffddc400007b56ffff84aaffffddc4;
    assign coff[1379] = 256'hffff909500003f01ffffc0ffffff909500006f6bffffc0ff00003f0100006f6b;
    assign coff[1380] = 256'h000060fdffffac7800005388000060fdffff9f0300005388ffffac78ffff9f03;
    assign coff[1381] = 256'hffff805bfffff67c00000984ffff805b00007fa500000984fffff67c00007fa5;
    assign coff[1382] = 256'hffffd7f1ffff866e00007992ffffd7f10000280f00007992ffff866e0000280f;
    assign coff[1383] = 256'hffffc65d0000724affff8db6ffffc65d000039a3ffff8db60000724a000039a3;
    assign coff[1384] = 256'h0000750fffffcc38000033c80000750fffff8af1000033c8ffffcc38ffff8af1;
    assign coff[1385] = 256'hffff889dffffd1d800002e28ffff889d0000776300002e28ffffd1d800007763;
    assign coff[1386] = 256'hfffffcf5ffff800900007ff7fffffcf50000030b00007ff7ffff80090000030b;
    assign coff[1387] = 256'hffffa7ab00005ca3ffffa35dffffa7ab00005855ffffa35d00005ca300005855;
    assign coff[1388] = 256'h00004490ffff93e900006c1700004490ffffbb7000006c17ffff93e9ffffbb70;
    assign coff[1389] = 256'hffff831700001bf3ffffe40dffff831700007ce9ffffe40d00001bf300007ce9;
    assign coff[1390] = 256'hffffb660ffff974b000068b5ffffb660000049a0000068b5ffff974b000049a0;
    assign coff[1391] = 256'hffffea0500007e19ffff81e7ffffea05000015fbffff81e700007e19000015fb;
    assign coff[1392] = 256'h00007b64ffffddf50000220b00007b64ffff849c0000220bffffddf5ffff849c;
    assign coff[1393] = 256'hffff90adffffc0d300003f2dffff90ad00006f5300003f2dffffc0d300006f53;
    assign coff[1394] = 256'h00000fc4ffff80fa00007f0600000fc4fffff03c00007f06ffff80fafffff03c;
    assign coff[1395] = 256'hffff9b0800004eacffffb154ffff9b08000064f8ffffb15400004eac000064f8;
    assign coff[1396] = 256'h000053aeffff9f24000060dc000053aeffffac52000060dcffff9f24ffffac52;
    assign coff[1397] = 256'hffff805700000951fffff6afffff805700007fa9fffff6af0000095100007fa9;
    assign coff[1398] = 256'hffffc68affff8da000007260ffffc68a0000397600007260ffff8da000003976;
    assign coff[1399] = 256'hffffd7c100007982ffff867effffd7c10000283fffff867e000079820000283f;
    assign coff[1400] = 256'h00006c32ffffbb9a0000446600006c32ffff93ce00004466ffffbb9affff93ce;
    assign coff[1401] = 256'hffff8322ffffe3dc00001c24ffff832200007cde00001c24ffffe3dc00007cde;
    assign coff[1402] = 256'hffffea37ffff81de00007e22ffffea37000015c900007e22ffff81de000015c9;
    assign coff[1403] = 256'hffffb63700006898ffff9768ffffb637000049c9ffff976800006898000049c9;
    assign coff[1404] = 256'h000033f6ffff8b05000074fb000033f6ffffcc0a000074fbffff8b05ffffcc0a;
    assign coff[1405] = 256'hffff888b00002dfaffffd206ffff888b00007775ffffd20600002dfa00007775;
    assign coff[1406] = 256'hffffa7cfffffa33b00005cc5ffffa7cf0000583100005cc5ffffa33b00005831;
    assign coff[1407] = 256'hfffffcc300007ff6ffff800afffffcc30000033dffff800a00007ff60000033d;
    assign coff[1408] = 256'h00007ff1fffffc2c000003d400007ff1ffff800f000003d4fffffc2cffff800f;
    assign coff[1409] = 256'hffffa2d3ffffa83d000057c3ffffa2d300005d2d000057c3ffffa83d00005d2d;
    assign coff[1410] = 256'h00002d6dffff8855000077ab00002d6dffffd293000077abffff8855ffffd293;
    assign coff[1411] = 256'hffff8b4300003480ffffcb80ffff8b43000074bdffffcb8000003480000074bd;
    assign coff[1412] = 256'h00006841ffffb5bc00004a4400006841ffff97bf00004a44ffffb5bcffff97bf;
    assign coff[1413] = 256'hffff81c5ffffeacb00001535ffff81c500007e3b00001535ffffeacb00007e3b;
    assign coff[1414] = 256'hffffe349ffff834300007cbdffffe34900001cb700007cbdffff834300001cb7;
    assign coff[1415] = 256'hffffbc1a00006c82ffff937effffbc1a000043e6ffff937e00006c82000043e6;
    assign coff[1416] = 256'h00007953ffffd732000028ce00007953ffff86ad000028ceffffd732ffff86ad;
    assign coff[1417] = 256'hffff8d5cffffc710000038f0ffff8d5c000072a4000038f0ffffc710000072a4;
    assign coff[1418] = 256'h000008bbffff804c00007fb4000008bbfffff74500007fb4ffff804cfffff745;
    assign coff[1419] = 256'hffff9f8700005420ffffabe0ffff9f8700006079ffffabe00000542000006079;
    assign coff[1420] = 256'h00004e35ffff9aac0000655400004e35ffffb1cb00006554ffff9aacffffb1cb;
    assign coff[1421] = 256'hffff810c0000105affffefa6ffff810c00007ef4ffffefa60000105a00007ef4;
    assign coff[1422] = 256'hffffc050ffff90f800006f08ffffc05000003fb000006f08ffff90f800003fb0;
    assign coff[1423] = 256'hffffde8600007b8bffff8475ffffde860000217affff847500007b8b0000217a;
    assign coff[1424] = 256'h00007dffffffe9710000168f00007dffffff82010000168fffffe971ffff8201;
    assign coff[1425] = 256'hffff96f4ffffb6dc00004924ffff96f40000690c00004924ffffb6dc0000690c;
    assign coff[1426] = 256'h00001b60ffff82f600007d0a00001b60ffffe4a000007d0affff82f6ffffe4a0;
    assign coff[1427] = 256'hffff943a0000450fffffbaf1ffff943a00006bc6ffffbaf10000450f00006bc6;
    assign coff[1428] = 256'h00005c3affffa73e000058c200005c3affffa3c6000058c2ffffa73effffa3c6;
    assign coff[1429] = 256'hffff8006fffffd8c00000274ffff800600007ffa00000274fffffd8c00007ffa;
    assign coff[1430] = 256'hffffd14bffff88d30000772dffffd14b00002eb50000772dffff88d300002eb5;
    assign coff[1431] = 256'hffffccc20000754cffff8ab4ffffccc20000333effff8ab40000754c0000333e;
    assign coff[1432] = 256'h00007206ffffc5d600003a2a00007206ffff8dfa00003a2affffc5d6ffff8dfa;
    assign coff[1433] = 256'hffff863fffffd88000002780ffff863f000079c100002780ffffd880000079c1;
    assign coff[1434] = 256'hfffff5e6ffff806600007f9afffff5e600000a1a00007f9affff806600000a1a;
    assign coff[1435] = 256'hffffacea0000615fffff9ea1ffffacea00005316ffff9ea10000615f00005316;
    assign coff[1436] = 256'h00003e7effff904b00006fb500003e7effffc18200006fb5ffff904bffffc182;
    assign coff[1437] = 256'hffff84d2000022cdffffdd33ffff84d200007b2effffdd33000022cd00007b2e;
    assign coff[1438] = 256'hffffb0b6ffff9b840000647cffffb0b600004f4a0000647cffff9b8400004f4a;
    assign coff[1439] = 256'hfffff10400007f1fffff80e1fffff10400000efcffff80e100007f1f00000efc;
    assign coff[1440] = 256'h00007f50fffff2c500000d3b00007f50ffff80b000000d3bfffff2c5ffff80b0;
    assign coff[1441] = 256'hffff9c9fffffaf54000050acffff9c9f00006361000050acffffaf5400006361;
    assign coff[1442] = 256'h00002480ffff855000007ab000002480ffffdb8000007ab0ffff8550ffffdb80;
    assign coff[1443] = 256'hffff8f7100003cf2ffffc30effff8f710000708fffffc30e00003cf20000708f;
    assign coff[1444] = 256'h00006282ffffae45000051bb00006282ffff9d7e000051bbffffae45ffff9d7e;
    assign coff[1445] = 256'hffff808dfffff42300000bddffff808d00007f7300000bddfffff42300007f73;
    assign coff[1446] = 256'hffffda30ffff85b700007a49ffffda30000025d000007a49ffff85b7000025d0;
    assign coff[1447] = 256'hffffc44500007135ffff8ecbffffc44500003bbbffff8ecb0000713500003bbb;
    assign coff[1448] = 256'h000075feffffce620000319e000075feffff8a020000319effffce62ffff8a02;
    assign coff[1449] = 256'hffff897bffffcfa700003059ffff897b0000768500003059ffffcfa700007685;
    assign coff[1450] = 256'hffffff50ffff800100007fffffffff50000000b000007fffffff8001000000b0;
    assign coff[1451] = 256'hffffa5fa00005affffffa501ffffa5fa00005a06ffffa50100005aff00005a06;
    assign coff[1452] = 256'h0000468affff953100006acf0000468affffb97600006acfffff9531ffffb976;
    assign coff[1453] = 256'hffff8298000019a5ffffe65bffff829800007d68ffffe65b000019a500007d68;
    assign coff[1454] = 256'hffffb851ffff95f500006a0bffffb851000047af00006a0bffff95f5000047af;
    assign coff[1455] = 256'hffffe7b400007dacffff8254ffffe7b40000184cffff825400007dac0000184c;
    assign coff[1456] = 256'h00007bffffffe03b00001fc500007bffffff840100001fc5ffffe03bffff8401;
    assign coff[1457] = 256'hffff91dcffffbec900004137ffff91dc00006e2400004137ffffbec900006e24;
    assign coff[1458] = 256'h0000121affff814900007eb70000121affffede600007eb7ffff8149ffffede6;
    assign coff[1459] = 256'hffff999a00004ccdffffb333ffff999a00006666ffffb33300004ccd00006666;
    assign coff[1460] = 256'h00005573ffffa0b300005f4d00005573ffffaa8d00005f4dffffa0b3ffffaa8d;
    assign coff[1461] = 256'hffff8031000006f8fffff908ffff803100007fcffffff908000006f800007fcf;
    assign coff[1462] = 256'hffffc8a7ffff8c960000736affffc8a7000037590000736affff8c9600003759;
    assign coff[1463] = 256'hffffd587000078bfffff8741ffffd58700002a79ffff8741000078bf00002a79;
    assign coff[1464] = 256'h00006d6fffffbd9b0000426500006d6fffff929100004265ffffbd9bffff9291;
    assign coff[1465] = 256'hffff83acffffe19100001e6fffff83ac00007c5400001e6fffffe19100007c54;
    assign coff[1466] = 256'hffffec8affff817d00007e83ffffec8a0000137600007e83ffff817d00001376;
    assign coff[1467] = 256'hffffb44e00006738ffff98c8ffffb44e00004bb2ffff98c80000673800004bb2;
    assign coff[1468] = 256'h0000361bffff8bff000074010000361bffffc9e500007401ffff8bffffffc9e5;
    assign coff[1469] = 256'hffff87b700002bc5ffffd43bffff87b700007849ffffd43b00002bc500007849;
    assign coff[1470] = 256'hffffa988ffffa19f00005e61ffffa9880000567800005e61ffffa19f00005678;
    assign coff[1471] = 256'hfffffa6800007fe1ffff801ffffffa6800000598ffff801f00007fe100000598;
    assign coff[1472] = 256'h00007fb7fffff7770000088900007fb7ffff804900000889fffff777ffff8049;
    assign coff[1473] = 256'hffff9fa8ffffabba00005446ffff9fa80000605800005446ffffabba00006058;
    assign coff[1474] = 256'h000028fdffff86be00007942000028fdffffd70300007942ffff86beffffd703;
    assign coff[1475] = 256'hffff8d46000038c2ffffc73effff8d46000072baffffc73e000038c2000072ba;
    assign coff[1476] = 256'h00006573ffffb1f300004e0d00006573ffff9a8d00004e0dffffb1f3ffff9a8d;
    assign coff[1477] = 256'hffff8113ffffef740000108cffff811300007eed0000108cffffef7400007eed;
    assign coff[1478] = 256'hffffdeb7ffff846700007b99ffffdeb70000214900007b99ffff846700002149;
    assign coff[1479] = 256'hffffc02400006eefffff9111ffffc02400003fdcffff911100006eef00003fdc;
    assign coff[1480] = 256'h000077bdffffd2c200002d3e000077bdffff884300002d3effffd2c2ffff8843;
    assign coff[1481] = 256'hffff8b58ffffcb53000034adffff8b58000074a8000034adffffcb53000074a8;
    assign coff[1482] = 256'h00000406ffff801000007ff000000406fffffbfa00007ff0ffff8010fffffbfa;
    assign coff[1483] = 256'hffffa2b00000579fffffa861ffffa2b000005d50ffffa8610000579f00005d50;
    assign coff[1484] = 256'h00004a6dffff97dc0000682400004a6dffffb59300006824ffff97dcffffb593;
    assign coff[1485] = 256'hffff81bd00001503ffffeafdffff81bd00007e43ffffeafd0000150300007e43;
    assign coff[1486] = 256'hffffbc45ffff936300006c9dffffbc45000043bb00006c9dffff9363000043bb;
    assign coff[1487] = 256'hffffe31800007cb1ffff834fffffe31800001ce8ffff834f00007cb100001ce8;
    assign coff[1488] = 256'h00007d15ffffe4d100001b2f00007d15ffff82eb00001b2fffffe4d1ffff82eb;
    assign coff[1489] = 256'hffff9456ffffbac700004539ffff945600006baa00004539ffffbac700006baa;
    assign coff[1490] = 256'h000016c1ffff820a00007df6000016c1ffffe93f00007df6ffff820affffe93f;
    assign coff[1491] = 256'hffff96d8000048fbffffb705ffff96d800006928ffffb705000048fb00006928;
    assign coff[1492] = 256'h000058e6ffffa3e800005c18000058e6ffffa71a00005c18ffffa3e8ffffa71a;
    assign coff[1493] = 256'hffff800500000242fffffdbeffff800500007ffbfffffdbe0000024200007ffb;
    assign coff[1494] = 256'hffffccf0ffff8aa000007560ffffccf00000331000007560ffff8aa000003310;
    assign coff[1495] = 256'hffffd11c0000771affff88e6ffffd11c00002ee4ffff88e60000771a00002ee4;
    assign coff[1496] = 256'h00006fceffffc1ae00003e5200006fceffff903200003e52ffffc1aeffff9032;
    assign coff[1497] = 256'hffff84e0ffffdd03000022fdffff84e000007b20000022fdffffdd0300007b20;
    assign coff[1498] = 256'hfffff135ffff80dc00007f24fffff13500000ecb00007f24ffff80dc00000ecb;
    assign coff[1499] = 256'hffffb08e0000645dffff9ba3ffffb08e00004f72ffff9ba30000645d00004f72;
    assign coff[1500] = 256'h00003a57ffff8e11000071ef00003a57ffffc5a9000071efffff8e11ffffc5a9;
    assign coff[1501] = 256'hffff863000002750ffffd8b0ffff8630000079d0ffffd8b000002750000079d0;
    assign coff[1502] = 256'hffffad11ffff9e810000617fffffad11000052ef0000617fffff9e81000052ef;
    assign coff[1503] = 256'hfffff5b400007f96ffff806afffff5b400000a4cffff806a00007f9600000a4c;
    assign coff[1504] = 256'h00007ebeffffee18000011e800007ebeffff8142000011e8ffffee18ffff8142;
    assign coff[1505] = 256'hffff99b8ffffb30b00004cf5ffff99b80000664800004cf5ffffb30b00006648;
    assign coff[1506] = 256'h00001ff5ffff840e00007bf200001ff5ffffe00b00007bf2ffff840effffe00b;
    assign coff[1507] = 256'hffff91c20000410cffffbef4ffff91c200006e3effffbef40000410c00006e3e;
    assign coff[1508] = 256'h00005f6fffffaab20000554e00005f6fffffa0910000554effffaab2ffffa091;
    assign coff[1509] = 256'hffff8033fffff8d60000072affff803300007fcd0000072afffff8d600007fcd;
    assign coff[1510] = 256'hffffd5b6ffff8730000078d0ffffd5b600002a4a000078d0ffff873000002a4a;
    assign coff[1511] = 256'hffffc87a00007355ffff8cabffffc87a00003786ffff8cab0000735500003786;
    assign coff[1512] = 256'h00007416ffffca13000035ed00007416ffff8bea000035edffffca13ffff8bea;
    assign coff[1513] = 256'hffff87c8ffffd40c00002bf4ffff87c80000783800002bf4ffffd40c00007838;
    assign coff[1514] = 256'hfffffa9affff801d00007fe3fffffa9a0000056600007fe3ffff801d00000566;
    assign coff[1515] = 256'hffffa96300005e3fffffa1c1ffffa9630000569dffffa1c100005e3f0000569d;
    assign coff[1516] = 256'h00004290ffff92ab00006d5500004290ffffbd7000006d55ffff92abffffbd70;
    assign coff[1517] = 256'hffff83a000001e3effffe1c2ffff83a000007c60ffffe1c200001e3e00007c60;
    assign coff[1518] = 256'hffffb476ffff98aa00006756ffffb47600004b8a00006756ffff98aa00004b8a;
    assign coff[1519] = 256'hffffec5800007e7bffff8185ffffec58000013a8ffff818500007e7b000013a8;
    assign coff[1520] = 256'h00007abeffffdbb10000244f00007abeffff85420000244fffffdbb1ffff8542;
    assign coff[1521] = 256'hffff8f89ffffc2e200003d1effff8f890000707700003d1effffc2e200007077;
    assign coff[1522] = 256'h00000d6dffff80b500007f4b00000d6dfffff29300007f4bffff80b5fffff293;
    assign coff[1523] = 256'hffff9c7f00005084ffffaf7cffff9c7f00006381ffffaf7c0000508400006381;
    assign coff[1524] = 256'h000051e2ffff9d9e00006262000051e2ffffae1e00006262ffff9d9effffae1e;
    assign coff[1525] = 256'hffff808800000babfffff455ffff808800007f78fffff45500000bab00007f78;
    assign coff[1526] = 256'hffffc471ffff8eb30000714dffffc47100003b8f0000714dffff8eb300003b8f;
    assign coff[1527] = 256'hffffda0000007a3bffff85c5ffffda0000002600ffff85c500007a3b00002600;
    assign coff[1528] = 256'h00006aebffffb9a00000466000006aebffff951500004660ffffb9a0ffff9515;
    assign coff[1529] = 256'hffff82a3ffffe62a000019d6ffff82a300007d5d000019d6ffffe62a00007d5d;
    assign coff[1530] = 256'hffffe7e5ffff824a00007db6ffffe7e50000181b00007db6ffff824a0000181b;
    assign coff[1531] = 256'hffffb827000069efffff9611ffffb827000047d9ffff9611000069ef000047d9;
    assign coff[1532] = 256'h000031ccffff8a16000075ea000031ccffffce34000075eaffff8a16ffffce34;
    assign coff[1533] = 256'hffff89680000302affffcfd6ffff896800007698ffffcfd60000302a00007698;
    assign coff[1534] = 256'hffffa61effffa4de00005b22ffffa61e000059e200005b22ffffa4de000059e2;
    assign coff[1535] = 256'hffffff1e00007fffffff8001ffffff1e000000e2ffff800100007fff000000e2;
    assign coff[1536] = 256'h00007fffffffff1e000000e200007fffffff8001000000e2ffffff1effff8001;
    assign coff[1537] = 256'hffffa4deffffa61e000059e2ffffa4de00005b22000059e2ffffa61e00005b22;
    assign coff[1538] = 256'h0000302affff8968000076980000302affffcfd600007698ffff8968ffffcfd6;
    assign coff[1539] = 256'hffff8a16000031ccffffce34ffff8a16000075eaffffce34000031cc000075ea;
    assign coff[1540] = 256'h000069efffffb827000047d9000069efffff9611000047d9ffffb827ffff9611;
    assign coff[1541] = 256'hffff824affffe7e50000181bffff824a00007db60000181bffffe7e500007db6;
    assign coff[1542] = 256'hffffe62affff82a300007d5dffffe62a000019d600007d5dffff82a3000019d6;
    assign coff[1543] = 256'hffffb9a000006aebffff9515ffffb9a000004660ffff951500006aeb00004660;
    assign coff[1544] = 256'h00007a3bffffda000000260000007a3bffff85c500002600ffffda00ffff85c5;
    assign coff[1545] = 256'hffff8eb3ffffc47100003b8fffff8eb30000714d00003b8fffffc4710000714d;
    assign coff[1546] = 256'h00000babffff808800007f7800000babfffff45500007f78ffff8088fffff455;
    assign coff[1547] = 256'hffff9d9e000051e2ffffae1effff9d9e00006262ffffae1e000051e200006262;
    assign coff[1548] = 256'h00005084ffff9c7f0000638100005084ffffaf7c00006381ffff9c7fffffaf7c;
    assign coff[1549] = 256'hffff80b500000d6dfffff293ffff80b500007f4bfffff29300000d6d00007f4b;
    assign coff[1550] = 256'hffffc2e2ffff8f8900007077ffffc2e200003d1e00007077ffff8f8900003d1e;
    assign coff[1551] = 256'hffffdbb100007abeffff8542ffffdbb10000244fffff854200007abe0000244f;
    assign coff[1552] = 256'h00007e7bffffec58000013a800007e7bffff8185000013a8ffffec58ffff8185;
    assign coff[1553] = 256'hffff98aaffffb47600004b8affff98aa0000675600004b8affffb47600006756;
    assign coff[1554] = 256'h00001e3effff83a000007c6000001e3effffe1c200007c60ffff83a0ffffe1c2;
    assign coff[1555] = 256'hffff92ab00004290ffffbd70ffff92ab00006d55ffffbd700000429000006d55;
    assign coff[1556] = 256'h00005e3fffffa9630000569d00005e3fffffa1c10000569dffffa963ffffa1c1;
    assign coff[1557] = 256'hffff801dfffffa9a00000566ffff801d00007fe300000566fffffa9a00007fe3;
    assign coff[1558] = 256'hffffd40cffff87c800007838ffffd40c00002bf400007838ffff87c800002bf4;
    assign coff[1559] = 256'hffffca1300007416ffff8beaffffca13000035edffff8bea00007416000035ed;
    assign coff[1560] = 256'h00007355ffffc87a0000378600007355ffff8cab00003786ffffc87affff8cab;
    assign coff[1561] = 256'hffff8730ffffd5b600002a4affff8730000078d000002a4affffd5b6000078d0;
    assign coff[1562] = 256'hfffff8d6ffff803300007fcdfffff8d60000072a00007fcdffff80330000072a;
    assign coff[1563] = 256'hffffaab200005f6fffffa091ffffaab20000554effffa09100005f6f0000554e;
    assign coff[1564] = 256'h0000410cffff91c200006e3e0000410cffffbef400006e3effff91c2ffffbef4;
    assign coff[1565] = 256'hffff840e00001ff5ffffe00bffff840e00007bf2ffffe00b00001ff500007bf2;
    assign coff[1566] = 256'hffffb30bffff99b800006648ffffb30b00004cf500006648ffff99b800004cf5;
    assign coff[1567] = 256'hffffee1800007ebeffff8142ffffee18000011e8ffff814200007ebe000011e8;
    assign coff[1568] = 256'h00007f96fffff5b400000a4c00007f96ffff806a00000a4cfffff5b4ffff806a;
    assign coff[1569] = 256'hffff9e81ffffad11000052efffff9e810000617f000052efffffad110000617f;
    assign coff[1570] = 256'h00002750ffff8630000079d000002750ffffd8b0000079d0ffff8630ffffd8b0;
    assign coff[1571] = 256'hffff8e1100003a57ffffc5a9ffff8e11000071efffffc5a900003a57000071ef;
    assign coff[1572] = 256'h0000645dffffb08e00004f720000645dffff9ba300004f72ffffb08effff9ba3;
    assign coff[1573] = 256'hffff80dcfffff13500000ecbffff80dc00007f2400000ecbfffff13500007f24;
    assign coff[1574] = 256'hffffdd03ffff84e000007b20ffffdd03000022fd00007b20ffff84e0000022fd;
    assign coff[1575] = 256'hffffc1ae00006fceffff9032ffffc1ae00003e52ffff903200006fce00003e52;
    assign coff[1576] = 256'h0000771affffd11c00002ee40000771affff88e600002ee4ffffd11cffff88e6;
    assign coff[1577] = 256'hffff8aa0ffffccf000003310ffff8aa00000756000003310ffffccf000007560;
    assign coff[1578] = 256'h00000242ffff800500007ffb00000242fffffdbe00007ffbffff8005fffffdbe;
    assign coff[1579] = 256'hffffa3e8000058e6ffffa71affffa3e800005c18ffffa71a000058e600005c18;
    assign coff[1580] = 256'h000048fbffff96d800006928000048fbffffb70500006928ffff96d8ffffb705;
    assign coff[1581] = 256'hffff820a000016c1ffffe93fffff820a00007df6ffffe93f000016c100007df6;
    assign coff[1582] = 256'hffffbac7ffff945600006baaffffbac70000453900006baaffff945600004539;
    assign coff[1583] = 256'hffffe4d100007d15ffff82ebffffe4d100001b2fffff82eb00007d1500001b2f;
    assign coff[1584] = 256'h00007cb1ffffe31800001ce800007cb1ffff834f00001ce8ffffe318ffff834f;
    assign coff[1585] = 256'hffff9363ffffbc45000043bbffff936300006c9d000043bbffffbc4500006c9d;
    assign coff[1586] = 256'h00001503ffff81bd00007e4300001503ffffeafd00007e43ffff81bdffffeafd;
    assign coff[1587] = 256'hffff97dc00004a6dffffb593ffff97dc00006824ffffb59300004a6d00006824;
    assign coff[1588] = 256'h0000579fffffa2b000005d500000579fffffa86100005d50ffffa2b0ffffa861;
    assign coff[1589] = 256'hffff801000000406fffffbfaffff801000007ff0fffffbfa0000040600007ff0;
    assign coff[1590] = 256'hffffcb53ffff8b58000074a8ffffcb53000034ad000074a8ffff8b58000034ad;
    assign coff[1591] = 256'hffffd2c2000077bdffff8843ffffd2c200002d3effff8843000077bd00002d3e;
    assign coff[1592] = 256'h00006eefffffc02400003fdc00006eefffff911100003fdcffffc024ffff9111;
    assign coff[1593] = 256'hffff8467ffffdeb700002149ffff846700007b9900002149ffffdeb700007b99;
    assign coff[1594] = 256'hffffef74ffff811300007eedffffef740000108c00007eedffff81130000108c;
    assign coff[1595] = 256'hffffb1f300006573ffff9a8dffffb1f300004e0dffff9a8d0000657300004e0d;
    assign coff[1596] = 256'h000038c2ffff8d46000072ba000038c2ffffc73e000072baffff8d46ffffc73e;
    assign coff[1597] = 256'hffff86be000028fdffffd703ffff86be00007942ffffd703000028fd00007942;
    assign coff[1598] = 256'hffffabbaffff9fa800006058ffffabba0000544600006058ffff9fa800005446;
    assign coff[1599] = 256'hfffff77700007fb7ffff8049fffff77700000889ffff804900007fb700000889;
    assign coff[1600] = 256'h00007fe1fffffa680000059800007fe1ffff801f00000598fffffa68ffff801f;
    assign coff[1601] = 256'hffffa19fffffa98800005678ffffa19f00005e6100005678ffffa98800005e61;
    assign coff[1602] = 256'h00002bc5ffff87b70000784900002bc5ffffd43b00007849ffff87b7ffffd43b;
    assign coff[1603] = 256'hffff8bff0000361bffffc9e5ffff8bff00007401ffffc9e50000361b00007401;
    assign coff[1604] = 256'h00006738ffffb44e00004bb200006738ffff98c800004bb2ffffb44effff98c8;
    assign coff[1605] = 256'hffff817dffffec8a00001376ffff817d00007e8300001376ffffec8a00007e83;
    assign coff[1606] = 256'hffffe191ffff83ac00007c54ffffe19100001e6f00007c54ffff83ac00001e6f;
    assign coff[1607] = 256'hffffbd9b00006d6fffff9291ffffbd9b00004265ffff929100006d6f00004265;
    assign coff[1608] = 256'h000078bfffffd58700002a79000078bfffff874100002a79ffffd587ffff8741;
    assign coff[1609] = 256'hffff8c96ffffc8a700003759ffff8c960000736a00003759ffffc8a70000736a;
    assign coff[1610] = 256'h000006f8ffff803100007fcf000006f8fffff90800007fcfffff8031fffff908;
    assign coff[1611] = 256'hffffa0b300005573ffffaa8dffffa0b300005f4dffffaa8d0000557300005f4d;
    assign coff[1612] = 256'h00004ccdffff999a0000666600004ccdffffb33300006666ffff999affffb333;
    assign coff[1613] = 256'hffff81490000121affffede6ffff814900007eb7ffffede60000121a00007eb7;
    assign coff[1614] = 256'hffffbec9ffff91dc00006e24ffffbec90000413700006e24ffff91dc00004137;
    assign coff[1615] = 256'hffffe03b00007bffffff8401ffffe03b00001fc5ffff840100007bff00001fc5;
    assign coff[1616] = 256'h00007dacffffe7b40000184c00007dacffff82540000184cffffe7b4ffff8254;
    assign coff[1617] = 256'hffff95f5ffffb851000047afffff95f500006a0b000047afffffb85100006a0b;
    assign coff[1618] = 256'h000019a5ffff829800007d68000019a5ffffe65b00007d68ffff8298ffffe65b;
    assign coff[1619] = 256'hffff95310000468affffb976ffff953100006acfffffb9760000468a00006acf;
    assign coff[1620] = 256'h00005affffffa5fa00005a0600005affffffa50100005a06ffffa5faffffa501;
    assign coff[1621] = 256'hffff8001ffffff50000000b0ffff800100007fff000000b0ffffff5000007fff;
    assign coff[1622] = 256'hffffcfa7ffff897b00007685ffffcfa70000305900007685ffff897b00003059;
    assign coff[1623] = 256'hffffce62000075feffff8a02ffffce620000319effff8a02000075fe0000319e;
    assign coff[1624] = 256'h00007135ffffc44500003bbb00007135ffff8ecb00003bbbffffc445ffff8ecb;
    assign coff[1625] = 256'hffff85b7ffffda30000025d0ffff85b700007a49000025d0ffffda3000007a49;
    assign coff[1626] = 256'hfffff423ffff808d00007f73fffff42300000bdd00007f73ffff808d00000bdd;
    assign coff[1627] = 256'hffffae4500006282ffff9d7effffae45000051bbffff9d7e00006282000051bb;
    assign coff[1628] = 256'h00003cf2ffff8f710000708f00003cf2ffffc30e0000708fffff8f71ffffc30e;
    assign coff[1629] = 256'hffff855000002480ffffdb80ffff855000007ab0ffffdb800000248000007ab0;
    assign coff[1630] = 256'hffffaf54ffff9c9f00006361ffffaf54000050ac00006361ffff9c9f000050ac;
    assign coff[1631] = 256'hfffff2c500007f50ffff80b0fffff2c500000d3bffff80b000007f5000000d3b;
    assign coff[1632] = 256'h00007f1ffffff10400000efc00007f1fffff80e100000efcfffff104ffff80e1;
    assign coff[1633] = 256'hffff9b84ffffb0b600004f4affff9b840000647c00004f4affffb0b60000647c;
    assign coff[1634] = 256'h000022cdffff84d200007b2e000022cdffffdd3300007b2effff84d2ffffdd33;
    assign coff[1635] = 256'hffff904b00003e7effffc182ffff904b00006fb5ffffc18200003e7e00006fb5;
    assign coff[1636] = 256'h0000615fffffacea000053160000615fffff9ea100005316ffffaceaffff9ea1;
    assign coff[1637] = 256'hffff8066fffff5e600000a1affff806600007f9a00000a1afffff5e600007f9a;
    assign coff[1638] = 256'hffffd880ffff863f000079c1ffffd88000002780000079c1ffff863f00002780;
    assign coff[1639] = 256'hffffc5d600007206ffff8dfaffffc5d600003a2affff8dfa0000720600003a2a;
    assign coff[1640] = 256'h0000754cffffccc20000333e0000754cffff8ab40000333effffccc2ffff8ab4;
    assign coff[1641] = 256'hffff88d3ffffd14b00002eb5ffff88d30000772d00002eb5ffffd14b0000772d;
    assign coff[1642] = 256'hfffffd8cffff800600007ffafffffd8c0000027400007ffaffff800600000274;
    assign coff[1643] = 256'hffffa73e00005c3affffa3c6ffffa73e000058c2ffffa3c600005c3a000058c2;
    assign coff[1644] = 256'h0000450fffff943a00006bc60000450fffffbaf100006bc6ffff943affffbaf1;
    assign coff[1645] = 256'hffff82f600001b60ffffe4a0ffff82f600007d0affffe4a000001b6000007d0a;
    assign coff[1646] = 256'hffffb6dcffff96f40000690cffffb6dc000049240000690cffff96f400004924;
    assign coff[1647] = 256'hffffe97100007dffffff8201ffffe9710000168fffff820100007dff0000168f;
    assign coff[1648] = 256'h00007b8bffffde860000217a00007b8bffff84750000217affffde86ffff8475;
    assign coff[1649] = 256'hffff90f8ffffc05000003fb0ffff90f800006f0800003fb0ffffc05000006f08;
    assign coff[1650] = 256'h0000105affff810c00007ef40000105affffefa600007ef4ffff810cffffefa6;
    assign coff[1651] = 256'hffff9aac00004e35ffffb1cbffff9aac00006554ffffb1cb00004e3500006554;
    assign coff[1652] = 256'h00005420ffff9f870000607900005420ffffabe000006079ffff9f87ffffabe0;
    assign coff[1653] = 256'hffff804c000008bbfffff745ffff804c00007fb4fffff745000008bb00007fb4;
    assign coff[1654] = 256'hffffc710ffff8d5c000072a4ffffc710000038f0000072a4ffff8d5c000038f0;
    assign coff[1655] = 256'hffffd73200007953ffff86adffffd732000028ceffff86ad00007953000028ce;
    assign coff[1656] = 256'h00006c82ffffbc1a000043e600006c82ffff937e000043e6ffffbc1affff937e;
    assign coff[1657] = 256'hffff8343ffffe34900001cb7ffff834300007cbd00001cb7ffffe34900007cbd;
    assign coff[1658] = 256'hffffeacbffff81c500007e3bffffeacb0000153500007e3bffff81c500001535;
    assign coff[1659] = 256'hffffb5bc00006841ffff97bfffffb5bc00004a44ffff97bf0000684100004a44;
    assign coff[1660] = 256'h00003480ffff8b43000074bd00003480ffffcb80000074bdffff8b43ffffcb80;
    assign coff[1661] = 256'hffff885500002d6dffffd293ffff8855000077abffffd29300002d6d000077ab;
    assign coff[1662] = 256'hffffa83dffffa2d300005d2dffffa83d000057c300005d2dffffa2d3000057c3;
    assign coff[1663] = 256'hfffffc2c00007ff1ffff800ffffffc2c000003d4ffff800f00007ff1000003d4;
    assign coff[1664] = 256'h00007ff6fffffcc30000033d00007ff6ffff800a0000033dfffffcc3ffff800a;
    assign coff[1665] = 256'hffffa33bffffa7cf00005831ffffa33b00005cc500005831ffffa7cf00005cc5;
    assign coff[1666] = 256'h00002dfaffff888b0000777500002dfaffffd20600007775ffff888bffffd206;
    assign coff[1667] = 256'hffff8b05000033f6ffffcc0affff8b05000074fbffffcc0a000033f6000074fb;
    assign coff[1668] = 256'h00006898ffffb637000049c900006898ffff9768000049c9ffffb637ffff9768;
    assign coff[1669] = 256'hffff81deffffea37000015c9ffff81de00007e22000015c9ffffea3700007e22;
    assign coff[1670] = 256'hffffe3dcffff832200007cdeffffe3dc00001c2400007cdeffff832200001c24;
    assign coff[1671] = 256'hffffbb9a00006c32ffff93ceffffbb9a00004466ffff93ce00006c3200004466;
    assign coff[1672] = 256'h00007982ffffd7c10000283f00007982ffff867e0000283fffffd7c1ffff867e;
    assign coff[1673] = 256'hffff8da0ffffc68a00003976ffff8da00000726000003976ffffc68a00007260;
    assign coff[1674] = 256'h00000951ffff805700007fa900000951fffff6af00007fa9ffff8057fffff6af;
    assign coff[1675] = 256'hffff9f24000053aeffffac52ffff9f24000060dcffffac52000053ae000060dc;
    assign coff[1676] = 256'h00004eacffff9b08000064f800004eacffffb154000064f8ffff9b08ffffb154;
    assign coff[1677] = 256'hffff80fa00000fc4fffff03cffff80fa00007f06fffff03c00000fc400007f06;
    assign coff[1678] = 256'hffffc0d3ffff90ad00006f53ffffc0d300003f2d00006f53ffff90ad00003f2d;
    assign coff[1679] = 256'hffffddf500007b64ffff849cffffddf50000220bffff849c00007b640000220b;
    assign coff[1680] = 256'h00007e19ffffea05000015fb00007e19ffff81e7000015fbffffea05ffff81e7;
    assign coff[1681] = 256'hffff974bffffb660000049a0ffff974b000068b5000049a0ffffb660000068b5;
    assign coff[1682] = 256'h00001bf3ffff831700007ce900001bf3ffffe40d00007ce9ffff8317ffffe40d;
    assign coff[1683] = 256'hffff93e900004490ffffbb70ffff93e900006c17ffffbb700000449000006c17;
    assign coff[1684] = 256'h00005ca3ffffa7ab0000585500005ca3ffffa35d00005855ffffa7abffffa35d;
    assign coff[1685] = 256'hffff8009fffffcf50000030bffff800900007ff70000030bfffffcf500007ff7;
    assign coff[1686] = 256'hffffd1d8ffff889d00007763ffffd1d800002e2800007763ffff889d00002e28;
    assign coff[1687] = 256'hffffcc380000750fffff8af1ffffcc38000033c8ffff8af10000750f000033c8;
    assign coff[1688] = 256'h0000724affffc65d000039a30000724affff8db6000039a3ffffc65dffff8db6;
    assign coff[1689] = 256'hffff866effffd7f10000280fffff866e000079920000280fffffd7f100007992;
    assign coff[1690] = 256'hfffff67cffff805b00007fa5fffff67c0000098400007fa5ffff805b00000984;
    assign coff[1691] = 256'hffffac78000060fdffff9f03ffffac7800005388ffff9f03000060fd00005388;
    assign coff[1692] = 256'h00003f01ffff909500006f6b00003f01ffffc0ff00006f6bffff9095ffffc0ff;
    assign coff[1693] = 256'hffff84aa0000223cffffddc4ffff84aa00007b56ffffddc40000223c00007b56;
    assign coff[1694] = 256'hffffb12cffff9b27000064d9ffffb12c00004ed4000064d9ffff9b2700004ed4;
    assign coff[1695] = 256'hfffff06e00007f0dffff80f3fffff06e00000f92ffff80f300007f0d00000f92;
    assign coff[1696] = 256'h00007f60fffff35b00000ca500007f60ffff80a000000ca5fffff35bffff80a0;
    assign coff[1697] = 256'hffff9cfeffffaee000005120ffff9cfe0000630200005120ffffaee000006302;
    assign coff[1698] = 256'h00002510ffff857c00007a8400002510ffffdaf000007a84ffff857cffffdaf0;
    assign coff[1699] = 256'hffff8f2900003c6dffffc393ffff8f29000070d7ffffc39300003c6d000070d7;
    assign coff[1700] = 256'h000062e2ffffaeb900005147000062e2ffff9d1e00005147ffffaeb9ffff9d1e;
    assign coff[1701] = 256'hffff809bfffff38d00000c73ffff809b00007f6500000c73fffff38d00007f65;
    assign coff[1702] = 256'hffffdac0ffff858a00007a76ffffdac00000254000007a76ffff858a00002540;
    assign coff[1703] = 256'hffffc3bf000070efffff8f11ffffc3bf00003c41ffff8f11000070ef00003c41;
    assign coff[1704] = 256'h00007638ffffceed0000311300007638ffff89c800003113ffffceedffff89c8;
    assign coff[1705] = 256'hffff89b5ffffcf1b000030e5ffff89b50000764b000030e5ffffcf1b0000764b;
    assign coff[1706] = 256'hffffffe7ffff800100007fffffffffe70000001900007fffffff800100000019;
    assign coff[1707] = 256'hffffa58f00005a94ffffa56cffffa58f00005a71ffffa56c00005a9400005a71;
    assign coff[1708] = 256'h00004708ffff958400006a7c00004708ffffb8f800006a7cffff9584ffffb8f8;
    assign coff[1709] = 256'hffff827b00001911ffffe6efffff827b00007d85ffffe6ef0000191100007d85;
    assign coff[1710] = 256'hffffb8ceffff95a000006a60ffffb8ce0000473200006a60ffff95a000004732;
    assign coff[1711] = 256'hffffe72000007d8fffff8271ffffe720000018e0ffff827100007d8f000018e0;
    assign coff[1712] = 256'h00007c24ffffe0ce00001f3200007c24ffff83dc00001f32ffffe0ceffff83dc;
    assign coff[1713] = 256'hffff9229ffffbe47000041b9ffff922900006dd7000041b9ffffbe4700006dd7;
    assign coff[1714] = 256'h000012afffff815f00007ea1000012afffffed5100007ea1ffff815fffffed51;
    assign coff[1715] = 256'hffff993f00004c54ffffb3acffff993f000066c1ffffb3ac00004c54000066c1;
    assign coff[1716] = 256'h000055e3ffffa11800005ee8000055e3ffffaa1d00005ee8ffffa118ffffaa1d;
    assign coff[1717] = 256'hffff802900000661fffff99fffff802900007fd7fffff99f0000066100007fd7;
    assign coff[1718] = 256'hffffc92fffff8c55000073abffffc92f000036d1000073abffff8c55000036d1;
    assign coff[1719] = 256'hffffd4f80000788dffff8773ffffd4f800002b08ffff87730000788d00002b08;
    assign coff[1720] = 256'h00006dbdffffbe1c000041e400006dbdffff9243000041e4ffffbe1cffff9243;
    assign coff[1721] = 256'hffff83d0ffffe0fe00001f02ffff83d000007c3000001f02ffffe0fe00007c30;
    assign coff[1722] = 256'hffffed1fffff816600007e9affffed1f000012e100007e9affff8166000012e1;
    assign coff[1723] = 256'hffffb3d4000066deffff9922ffffb3d400004c2cffff9922000066de00004c2c;
    assign coff[1724] = 256'h000036a3ffff8c3f000073c1000036a3ffffc95d000073c1ffff8c3fffffc95d;
    assign coff[1725] = 256'hffff878400002b37ffffd4c9ffff87840000787cffffd4c900002b370000787c;
    assign coff[1726] = 256'hffffa9f8ffffa13900005ec7ffffa9f80000560800005ec7ffffa13900005608;
    assign coff[1727] = 256'hfffff9d100007fdaffff8026fffff9d10000062fffff802600007fda0000062f;
    assign coff[1728] = 256'h00007fc1fffff80e000007f200007fc1ffff803f000007f2fffff80effff803f;
    assign coff[1729] = 256'hffffa00cffffab49000054b7ffffa00c00005ff4000054b7ffffab4900005ff4;
    assign coff[1730] = 256'h0000298cffff86ee000079120000298cffffd67400007912ffff86eeffffd674;
    assign coff[1731] = 256'hffff8d030000383bffffc7c5ffff8d03000072fdffffc7c50000383b000072fd;
    assign coff[1732] = 256'h000065cfffffb26b00004d95000065cfffff9a3100004d95ffffb26bffff9a31;
    assign coff[1733] = 256'hffff8127ffffeedf00001121ffff812700007ed900001121ffffeedf00007ed9;
    assign coff[1734] = 256'hffffdf48ffff844100007bbfffffdf48000020b800007bbfffff8441000020b8;
    assign coff[1735] = 256'hffffbfa200006ea3ffff915dffffbfa20000405effff915d00006ea30000405e;
    assign coff[1736] = 256'h000077f2ffffd34f00002cb1000077f2ffff880e00002cb1ffffd34fffff880e;
    assign coff[1737] = 256'hffff8b96ffffcac900003537ffff8b960000746a00003537ffffcac90000746a;
    assign coff[1738] = 256'h0000049dffff801500007feb0000049dfffffb6300007febffff8015fffffb63;
    assign coff[1739] = 256'hffffa24900005730ffffa8d0ffffa24900005db7ffffa8d00000573000005db7;
    assign coff[1740] = 256'h00004ae7ffff9834000067cc00004ae7ffffb519000067ccffff9834ffffb519;
    assign coff[1741] = 256'hffff81a40000146effffeb92ffff81a400007e5cffffeb920000146e00007e5c;
    assign coff[1742] = 256'hffffbcc5ffff931400006cecffffbcc50000433b00006cecffff93140000433b;
    assign coff[1743] = 256'hffffe28500007c8fffff8371ffffe28500001d7bffff837100007c8f00001d7b;
    assign coff[1744] = 256'h00007d34ffffe56500001a9b00007d34ffff82cc00001a9bffffe565ffff82cc;
    assign coff[1745] = 256'hffff94a7ffffba48000045b8ffff94a700006b59000045b8ffffba4800006b59;
    assign coff[1746] = 256'h00001755ffff822500007ddb00001755ffffe8ab00007ddbffff8225ffffe8ab;
    assign coff[1747] = 256'hffff96820000487fffffb781ffff96820000697effffb7810000487f0000697e;
    assign coff[1748] = 256'h00005952ffffa45100005baf00005952ffffa6ae00005bafffffa451ffffa6ae;
    assign coff[1749] = 256'hffff8003000001abfffffe55ffff800300007ffdfffffe55000001ab00007ffd;
    assign coff[1750] = 256'hffffcd7bffff8a640000759cffffcd7b000032850000759cffff8a6400003285;
    assign coff[1751] = 256'hffffd090000076e3ffff891dffffd09000002f70ffff891d000076e300002f70;
    assign coff[1752] = 256'h00007017ffffc23200003dce00007017ffff8fe900003dceffffc232ffff8fe9;
    assign coff[1753] = 256'hffff850affffdc720000238effff850a00007af60000238effffdc7200007af6;
    assign coff[1754] = 256'hfffff1cbffff80ca00007f36fffff1cb00000e3500007f36ffff80ca00000e35;
    assign coff[1755] = 256'hffffb018000063ffffff9c01ffffb01800004fe8ffff9c01000063ff00004fe8;
    assign coff[1756] = 256'h00003addffff8e56000071aa00003addffffc523000071aaffff8e56ffffc523;
    assign coff[1757] = 256'hffff8602000026c0ffffd940ffff8602000079feffffd940000026c0000079fe;
    assign coff[1758] = 256'hffffad84ffff9e1f000061e1ffffad840000527c000061e1ffff9e1f0000527c;
    assign coff[1759] = 256'hfffff51e00007f89ffff8077fffff51e00000ae2ffff807700007f8900000ae2;
    assign coff[1760] = 256'h00007ed3ffffeead0000115300007ed3ffff812d00001153ffffeeadffff812d;
    assign coff[1761] = 256'hffff9a13ffffb29300004d6dffff9a13000065ed00004d6dffffb293000065ed;
    assign coff[1762] = 256'h00002087ffff843400007bcc00002087ffffdf7900007bccffff8434ffffdf79;
    assign coff[1763] = 256'hffff91760000408affffbf76ffff917600006e8affffbf760000408a00006e8a;
    assign coff[1764] = 256'h00005fd3ffffab23000054dd00005fd3ffffa02d000054ddffffab23ffffa02d;
    assign coff[1765] = 256'hffff803cfffff840000007c0ffff803c00007fc4000007c0fffff84000007fc4;
    assign coff[1766] = 256'hffffd644ffff86ff00007901ffffd644000029bc00007901ffff86ff000029bc;
    assign coff[1767] = 256'hffffc7f200007313ffff8cedffffc7f20000380effff8ced000073130000380e;
    assign coff[1768] = 256'h00007455ffffca9c0000356400007455ffff8bab00003564ffffca9cffff8bab;
    assign coff[1769] = 256'hffff87fdffffd37f00002c81ffff87fd0000780300002c81ffffd37f00007803;
    assign coff[1770] = 256'hfffffb31ffff801700007fe9fffffb31000004cf00007fe9ffff8017000004cf;
    assign coff[1771] = 256'hffffa8f400005dd9ffffa227ffffa8f40000570cffffa22700005dd90000570c;
    assign coff[1772] = 256'h00004310ffff92fa00006d0600004310ffffbcf000006d06ffff92faffffbcf0;
    assign coff[1773] = 256'hffff837d00001dacffffe254ffff837d00007c83ffffe25400001dac00007c83;
    assign coff[1774] = 256'hffffb4f0ffff9852000067aeffffb4f000004b10000067aeffff985200004b10;
    assign coff[1775] = 256'hffffebc300007e64ffff819cffffebc30000143dffff819c00007e640000143d;
    assign coff[1776] = 256'h00007ae8ffffdc41000023bf00007ae8ffff8518000023bfffffdc41ffff8518;
    assign coff[1777] = 256'hffff8fd1ffffc25e00003da2ffff8fd10000702f00003da2ffffc25e0000702f;
    assign coff[1778] = 256'h00000e03ffff80c500007f3b00000e03fffff1fd00007f3bffff80c5fffff1fd;
    assign coff[1779] = 256'hffff9c210000500fffffaff1ffff9c21000063dfffffaff10000500f000063df;
    assign coff[1780] = 256'h00005256ffff9dff0000620100005256ffffadaa00006201ffff9dffffffadaa;
    assign coff[1781] = 256'hffff807b00000b14fffff4ecffff807b00007f85fffff4ec00000b1400007f85;
    assign coff[1782] = 256'hffffc4f7ffff8e6d00007193ffffc4f700003b0900007193ffff8e6d00003b09;
    assign coff[1783] = 256'hffffd97000007a0effff85f2ffffd97000002690ffff85f200007a0e00002690;
    assign coff[1784] = 256'h00006b3dffffba1e000045e200006b3dffff94c3000045e2ffffba1effff94c3;
    assign coff[1785] = 256'hffff82c1ffffe59600001a6affff82c100007d3f00001a6affffe59600007d3f;
    assign coff[1786] = 256'hffffe879ffff822e00007dd2ffffe8790000178700007dd2ffff822e00001787;
    assign coff[1787] = 256'hffffb7ab0000699affff9666ffffb7ab00004855ffff96660000699a00004855;
    assign coff[1788] = 256'h00003257ffff8a51000075af00003257ffffcda9000075afffff8a51ffffcda9;
    assign coff[1789] = 256'hffff893000002f9fffffd061ffff8930000076d0ffffd06100002f9f000076d0;
    assign coff[1790] = 256'hffffa68affffa47400005b8cffffa68a0000597600005b8cffffa47400005976;
    assign coff[1791] = 256'hfffffe8700007ffeffff8002fffffe8700000179ffff800200007ffe00000179;
    assign coff[1792] = 256'h00007ffcfffffdf00000021000007ffcffff800400000210fffffdf0ffff8004;
    assign coff[1793] = 256'hffffa40bffffa6f60000590affffa40b00005bf50000590affffa6f600005bf5;
    assign coff[1794] = 256'h00002f13ffff88f80000770800002f13ffffd0ed00007708ffff88f8ffffd0ed;
    assign coff[1795] = 256'hffff8a8c000032e2ffffcd1effff8a8c00007574ffffcd1e000032e200007574;
    assign coff[1796] = 256'h00006945ffffb72f000048d100006945ffff96bb000048d1ffffb72fffff96bb;
    assign coff[1797] = 256'hffff8213ffffe90e000016f2ffff821300007ded000016f2ffffe90e00007ded;
    assign coff[1798] = 256'hffffe502ffff82e100007d1fffffe50200001afe00007d1fffff82e100001afe;
    assign coff[1799] = 256'hffffba9c00006b8fffff9471ffffba9c00004564ffff947100006b8f00004564;
    assign coff[1800] = 256'h000079e0ffffd8e000002720000079e0ffff862000002720ffffd8e0ffff8620;
    assign coff[1801] = 256'hffff8e28ffffc57d00003a83ffff8e28000071d800003a83ffffc57d000071d8;
    assign coff[1802] = 256'h00000a7effff806e00007f9200000a7efffff58200007f92ffff806efffff582;
    assign coff[1803] = 256'hffff9e60000052c9ffffad37ffff9e60000061a0ffffad37000052c9000061a0;
    assign coff[1804] = 256'h00004f99ffff9bc20000643e00004f99ffffb0670000643effff9bc2ffffb067;
    assign coff[1805] = 256'hffff80d600000e99fffff167ffff80d600007f2afffff16700000e9900007f2a;
    assign coff[1806] = 256'hffffc1daffff901a00006fe6ffffc1da00003e2600006fe6ffff901a00003e26;
    assign coff[1807] = 256'hffffdcd200007b12ffff84eeffffdcd20000232effff84ee00007b120000232e;
    assign coff[1808] = 256'h00007e4cffffeb2f000014d100007e4cffff81b4000014d1ffffeb2fffff81b4;
    assign coff[1809] = 256'hffff97faffffb56b00004a95ffff97fa0000680600004a95ffffb56b00006806;
    assign coff[1810] = 256'h00001d19ffff835a00007ca600001d19ffffe2e700007ca6ffff835affffe2e7;
    assign coff[1811] = 256'hffff934900004391ffffbc6fffff934900006cb7ffffbc6f0000439100006cb7;
    assign coff[1812] = 256'h00005d72ffffa8860000577a00005d72ffffa28e0000577affffa886ffffa28e;
    assign coff[1813] = 256'hffff8012fffffbc700000439ffff801200007fee00000439fffffbc700007fee;
    assign coff[1814] = 256'hffffd2f1ffff8831000077cfffffd2f100002d0f000077cfffff883100002d0f;
    assign coff[1815] = 256'hffffcb2500007494ffff8b6cffffcb25000034dbffff8b6c00007494000034db;
    assign coff[1816] = 256'h000072d0ffffc76b00003895000072d0ffff8d3000003895ffffc76bffff8d30;
    assign coff[1817] = 256'hffff86ceffffd6d30000292dffff86ce000079320000292dffffd6d300007932;
    assign coff[1818] = 256'hfffff7a9ffff804600007fbafffff7a90000085700007fbaffff804600000857;
    assign coff[1819] = 256'hffffab9400006037ffff9fc9ffffab940000546cffff9fc9000060370000546c;
    assign coff[1820] = 256'h00004007ffff912a00006ed600004007ffffbff900006ed6ffff912affffbff9;
    assign coff[1821] = 256'hffff845a00002119ffffdee7ffff845a00007ba6ffffdee70000211900007ba6;
    assign coff[1822] = 256'hffffb21bffff9a6e00006592ffffb21b00004de500006592ffff9a6e00004de5;
    assign coff[1823] = 256'hffffef4300007ee7ffff8119ffffef43000010bdffff811900007ee7000010bd;
    assign coff[1824] = 256'h00007f7cfffff48700000b7900007f7cffff808400000b79fffff487ffff8084;
    assign coff[1825] = 256'hffff9dbeffffadf700005209ffff9dbe0000624200005209ffffadf700006242;
    assign coff[1826] = 256'h00002630ffff85d400007a2c00002630ffffd9d000007a2cffff85d4ffffd9d0;
    assign coff[1827] = 256'hffff8e9c00003b62ffffc49effff8e9c00007164ffffc49e00003b6200007164;
    assign coff[1828] = 256'h000063a0ffffafa30000505d000063a0ffff9c600000505dffffafa3ffff9c60;
    assign coff[1829] = 256'hffff80bafffff26100000d9fffff80ba00007f4600000d9ffffff26100007f46;
    assign coff[1830] = 256'hffffdbe1ffff853400007accffffdbe10000241f00007accffff85340000241f;
    assign coff[1831] = 256'hffffc2b60000705fffff8fa1ffffc2b600003d4affff8fa10000705f00003d4a;
    assign coff[1832] = 256'h000076aaffffd00400002ffc000076aaffff895600002ffcffffd004ffff8956;
    assign coff[1833] = 256'hffff8a29ffffce05000031fbffff8a29000075d7000031fbffffce05000075d7;
    assign coff[1834] = 256'h00000114ffff800100007fff00000114fffffeec00007fffffff8001fffffeec;
    assign coff[1835] = 256'hffffa4bb000059beffffa642ffffa4bb00005b45ffffa642000059be00005b45;
    assign coff[1836] = 256'h00004802ffff962d000069d300004802ffffb7fe000069d3ffff962dffffb7fe;
    assign coff[1837] = 256'hffff8241000017e9ffffe817ffff824100007dbfffffe817000017e900007dbf;
    assign coff[1838] = 256'hffffb9caffff94fa00006b06ffffb9ca0000463600006b06ffff94fa00004636;
    assign coff[1839] = 256'hffffe5f800007d53ffff82adffffe5f800001a08ffff82ad00007d5300001a08;
    assign coff[1840] = 256'h00007c6cffffe1f200001e0e00007c6cffff839400001e0effffe1f2ffff8394;
    assign coff[1841] = 256'hffff92c5ffffbd45000042bbffff92c500006d3b000042bbffffbd4500006d3b;
    assign coff[1842] = 256'h000013d9ffff818c00007e74000013d9ffffec2700007e74ffff818cffffec27;
    assign coff[1843] = 256'hffff988d00004b61ffffb49fffff988d00006773ffffb49f00004b6100006773;
    assign coff[1844] = 256'h000056c2ffffa1e300005e1d000056c2ffffa93e00005e1dffffa1e3ffffa93e;
    assign coff[1845] = 256'hffff801b00000534fffffaccffff801b00007fe5fffffacc0000053400007fe5;
    assign coff[1846] = 256'hffffca40ffff8bd50000742bffffca40000035c00000742bffff8bd5000035c0;
    assign coff[1847] = 256'hffffd3dd00007826ffff87daffffd3dd00002c23ffff87da0000782600002c23;
    assign coff[1848] = 256'h00006e57ffffbf20000040e000006e57ffff91a9000040e0ffffbf20ffff91a9;
    assign coff[1849] = 256'hffff841affffdfda00002026ffff841a00007be600002026ffffdfda00007be6;
    assign coff[1850] = 256'hffffee4affff813b00007ec5ffffee4a000011b600007ec5ffff813b000011b6;
    assign coff[1851] = 256'hffffb2e30000662affff99d6ffffb2e300004d1dffff99d60000662a00004d1d;
    assign coff[1852] = 256'h000037b4ffff8cc10000733f000037b4ffffc84c0000733fffff8cc1ffffc84c;
    assign coff[1853] = 256'hffff871f00002a1bffffd5e5ffff871f000078e1ffffd5e500002a1b000078e1;
    assign coff[1854] = 256'hffffaad8ffffa07000005f90ffffaad80000552800005f90ffffa07000005528;
    assign coff[1855] = 256'hfffff8a400007fcaffff8036fffff8a40000075cffff803600007fca0000075c;
    assign coff[1856] = 256'h00007fd2fffff93b000006c500007fd2ffff802e000006c5fffff93bffff802e;
    assign coff[1857] = 256'hffffa0d4ffffaa6800005598ffffa0d400005f2c00005598ffffaa6800005f2c;
    assign coff[1858] = 256'h00002aa9ffff8751000078af00002aa9ffffd557000078afffff8751ffffd557;
    assign coff[1859] = 256'hffff8c800000372cffffc8d4ffff8c8000007380ffffc8d40000372c00007380;
    assign coff[1860] = 256'h00006684ffffb35b00004ca500006684ffff997c00004ca5ffffb35bffff997c;
    assign coff[1861] = 256'hffff8150ffffedb40000124cffff815000007eb00000124cffffedb400007eb0;
    assign coff[1862] = 256'hffffe06cffff83f500007c0bffffe06c00001f9400007c0bffff83f500001f94;
    assign coff[1863] = 256'hffffbe9e00006e0affff91f6ffffbe9e00004162ffff91f600006e0a00004162;
    assign coff[1864] = 256'h0000785affffd46b00002b950000785affff87a600002b95ffffd46bffff87a6;
    assign coff[1865] = 256'hffff8c15ffffc9b800003648ffff8c15000073eb00003648ffffc9b8000073eb;
    assign coff[1866] = 256'h000005caffff802200007fde000005cafffffa3600007fdeffff8022fffffa36;
    assign coff[1867] = 256'hffffa17d00005653ffffa9adffffa17d00005e83ffffa9ad0000565300005e83;
    assign coff[1868] = 256'h00004bdbffff98e60000671a00004bdbffffb4250000671affff98e6ffffb425;
    assign coff[1869] = 256'hffff817500001344ffffecbcffff817500007e8bffffecbc0000134400007e8b;
    assign coff[1870] = 256'hffffbdc6ffff927700006d89ffffbdc60000423a00006d89ffff92770000423a;
    assign coff[1871] = 256'hffffe16000007c48ffff83b8ffffe16000001ea0ffff83b800007c4800001ea0;
    assign coff[1872] = 256'h00007d72ffffe68c0000197400007d72ffff828e00001974ffffe68cffff828e;
    assign coff[1873] = 256'hffff954dffffb94c000046b4ffff954d00006ab3000046b4ffffb94c00006ab3;
    assign coff[1874] = 256'h0000187dffff825d00007da30000187dffffe78300007da3ffff825dffffe783;
    assign coff[1875] = 256'hffff95d800004785ffffb87bffff95d800006a28ffffb87b0000478500006a28;
    assign coff[1876] = 256'h00005a29ffffa52500005adb00005a29ffffa5d700005adbffffa525ffffa5d7;
    assign coff[1877] = 256'hffff80010000007effffff82ffff800100007fffffffff820000007e00007fff;
    assign coff[1878] = 256'hffffce90ffff89ef00007611ffffce900000317000007611ffff89ef00003170;
    assign coff[1879] = 256'hffffcf7800007672ffff898effffcf7800003088ffff898e0000767200003088;
    assign coff[1880] = 256'h000070a7ffffc33b00003cc5000070a7ffff8f5900003cc5ffffc33bffff8f59;
    assign coff[1881] = 256'hffff855fffffdb50000024b0ffff855f00007aa1000024b0ffffdb5000007aa1;
    assign coff[1882] = 256'hfffff2f7ffff80aa00007f56fffff2f700000d0900007f56ffff80aa00000d09;
    assign coff[1883] = 256'hffffaf2d00006342ffff9cbeffffaf2d000050d3ffff9cbe00006342000050d3;
    assign coff[1884] = 256'h00003be8ffff8ee20000711e00003be8ffffc4180000711effff8ee2ffffc418;
    assign coff[1885] = 256'hffff85a8000025a0ffffda60ffff85a800007a58ffffda60000025a000007a58;
    assign coff[1886] = 256'hffffae6bffff9d5e000062a2ffffae6b00005195000062a2ffff9d5e00005195;
    assign coff[1887] = 256'hfffff3f100007f6effff8092fffff3f100000c0fffff809200007f6e00000c0f;
    assign coff[1888] = 256'h00007efaffffefd80000102800007efaffff810600001028ffffefd8ffff8106;
    assign coff[1889] = 256'hffff9acaffffb1a300004e5dffff9aca0000653600004e5dffffb1a300006536;
    assign coff[1890] = 256'h000021aaffff848200007b7e000021aaffffde5600007b7effff8482ffffde56;
    assign coff[1891] = 256'hffff90df00003f85ffffc07bffff90df00006f21ffffc07b00003f8500006f21;
    assign coff[1892] = 256'h0000609affffac06000053fa0000609affff9f66000053faffffac06ffff9f66;
    assign coff[1893] = 256'hffff8050fffff713000008edffff805000007fb0000008edfffff71300007fb0;
    assign coff[1894] = 256'hffffd762ffff869e00007962ffffd7620000289e00007962ffff869e0000289e;
    assign coff[1895] = 256'hffffc6e30000728dffff8d73ffffc6e30000391dffff8d730000728d0000391d;
    assign coff[1896] = 256'h000074d2ffffcbae00003452000074d2ffff8b2e00003452ffffcbaeffff8b2e;
    assign coff[1897] = 256'hffff8867ffffd26400002d9cffff88670000779900002d9cffffd26400007799;
    assign coff[1898] = 256'hfffffc5effff800d00007ff3fffffc5e000003a200007ff3ffff800d000003a2;
    assign coff[1899] = 256'hffffa81800005d0bffffa2f5ffffa818000057e8ffffa2f500005d0b000057e8;
    assign coff[1900] = 256'h00004411ffff939900006c6700004411ffffbbef00006c67ffff9399ffffbbef;
    assign coff[1901] = 256'hffff833800001c86ffffe37affff833800007cc8ffffe37a00001c8600007cc8;
    assign coff[1902] = 256'hffffb5e5ffff97a20000685effffb5e500004a1b0000685effff97a200004a1b;
    assign coff[1903] = 256'hffffea9a00007e33ffff81cdffffea9a00001566ffff81cd00007e3300001566;
    assign coff[1904] = 256'h00007b3bffffdd630000229d00007b3bffff84c50000229dffffdd63ffff84c5;
    assign coff[1905] = 256'hffff9063ffffc15600003eaaffff906300006f9d00003eaaffffc15600006f9d;
    assign coff[1906] = 256'h00000f2effff80e700007f1900000f2efffff0d200007f19ffff80e7fffff0d2;
    assign coff[1907] = 256'hffff9b6500004f23ffffb0ddffff9b650000649bffffb0dd00004f230000649b;
    assign coff[1908] = 256'h0000533cffff9ec20000613e0000533cffffacc40000613effff9ec2ffffacc4;
    assign coff[1909] = 256'hffff8062000009e8fffff618ffff806200007f9efffff618000009e800007f9e;
    assign coff[1910] = 256'hffffc603ffff8de40000721cffffc603000039fd0000721cffff8de4000039fd;
    assign coff[1911] = 256'hffffd851000079b1ffff864fffffd851000027afffff864f000079b1000027af;
    assign coff[1912] = 256'h00006be1ffffbb1b000044e500006be1ffff941f000044e5ffffbb1bffff941f;
    assign coff[1913] = 256'hffff8301ffffe46f00001b91ffff830100007cff00001b91ffffe46f00007cff;
    assign coff[1914] = 256'hffffe9a2ffff81f800007e08ffffe9a20000165e00007e08ffff81f80000165e;
    assign coff[1915] = 256'hffffb6b3000068efffff9711ffffb6b30000494dffff9711000068ef0000494d;
    assign coff[1916] = 256'h0000336cffff8ac8000075380000336cffffcc9400007538ffff8ac8ffffcc94;
    assign coff[1917] = 256'hffff88c100002e86ffffd17affff88c10000773fffffd17a00002e860000773f;
    assign coff[1918] = 256'hffffa762ffffa3a300005c5dffffa7620000589e00005c5dffffa3a30000589e;
    assign coff[1919] = 256'hfffffd5900007ff9ffff8007fffffd59000002a7ffff800700007ff9000002a7;
    assign coff[1920] = 256'h00007fecfffffb950000046b00007fecffff80140000046bfffffb95ffff8014;
    assign coff[1921] = 256'hffffa26cffffa8ab00005755ffffa26c00005d9400005755ffffa8ab00005d94;
    assign coff[1922] = 256'h00002ce0ffff8820000077e000002ce0ffffd320000077e0ffff8820ffffd320;
    assign coff[1923] = 256'hffff8b8100003509ffffcaf7ffff8b810000747fffffcaf7000035090000747f;
    assign coff[1924] = 256'h000067e9ffffb54200004abe000067e9ffff981700004abeffffb542ffff9817;
    assign coff[1925] = 256'hffff81acffffeb60000014a0ffff81ac00007e54000014a0ffffeb6000007e54;
    assign coff[1926] = 256'hffffe2b6ffff836500007c9bffffe2b600001d4a00007c9bffff836500001d4a;
    assign coff[1927] = 256'hffffbc9a00006cd2ffff932effffbc9a00004366ffff932e00006cd200004366;
    assign coff[1928] = 256'h00007922ffffd6a40000295c00007922ffff86de0000295cffffd6a4ffff86de;
    assign coff[1929] = 256'hffff8d19ffffc79800003868ffff8d19000072e700003868ffffc798000072e7;
    assign coff[1930] = 256'h00000825ffff804200007fbe00000825fffff7db00007fbeffff8042fffff7db;
    assign coff[1931] = 256'hffff9fea00005491ffffab6fffff9fea00006016ffffab6f0000549100006016;
    assign coff[1932] = 256'h00004dbdffff9a50000065b000004dbdffffb243000065b0ffff9a50ffffb243;
    assign coff[1933] = 256'hffff8120000010efffffef11ffff812000007ee0ffffef11000010ef00007ee0;
    assign coff[1934] = 256'hffffbfcdffff914300006ebdffffbfcd0000403300006ebdffff914300004033;
    assign coff[1935] = 256'hffffdf1800007bb3ffff844dffffdf18000020e8ffff844d00007bb3000020e8;
    assign coff[1936] = 256'h00007de4ffffe8dc0000172400007de4ffff821c00001724ffffe8dcffff821c;
    assign coff[1937] = 256'hffff969fffffb758000048a8ffff969f00006961000048a8ffffb75800006961;
    assign coff[1938] = 256'h00001accffff82d600007d2a00001accffffe53400007d2affff82d6ffffe534;
    assign coff[1939] = 256'hffff948c0000458effffba72ffff948c00006b74ffffba720000458e00006b74;
    assign coff[1940] = 256'h00005bd2ffffa6d20000592e00005bd2ffffa42e0000592effffa6d2ffffa42e;
    assign coff[1941] = 256'hffff8003fffffe22000001deffff800300007ffd000001defffffe2200007ffd;
    assign coff[1942] = 256'hffffd0bfffff890b000076f5ffffd0bf00002f41000076f5ffff890b00002f41;
    assign coff[1943] = 256'hffffcd4c00007588ffff8a78ffffcd4c000032b4ffff8a7800007588000032b4;
    assign coff[1944] = 256'h000071c1ffffc55000003ab0000071c1ffff8e3f00003ab0ffffc550ffff8e3f;
    assign coff[1945] = 256'hffff8611ffffd910000026f0ffff8611000079ef000026f0ffffd910000079ef;
    assign coff[1946] = 256'hfffff550ffff807200007f8efffff55000000ab000007f8effff807200000ab0;
    assign coff[1947] = 256'hffffad5d000061c0ffff9e40ffffad5d000052a3ffff9e40000061c0000052a3;
    assign coff[1948] = 256'h00003dfaffff900100006fff00003dfaffffc20600006fffffff9001ffffc206;
    assign coff[1949] = 256'hffff84fc0000235effffdca2ffff84fc00007b04ffffdca20000235e00007b04;
    assign coff[1950] = 256'hffffb040ffff9be20000641effffb04000004fc00000641effff9be200004fc0;
    assign coff[1951] = 256'hfffff19900007f30ffff80d0fffff19900000e67ffff80d000007f3000000e67;
    assign coff[1952] = 256'h00007f41fffff22f00000dd100007f41ffff80bf00000dd1fffff22fffff80bf;
    assign coff[1953] = 256'hffff9c40ffffafca00005036ffff9c40000063c000005036ffffafca000063c0;
    assign coff[1954] = 256'h000023efffff852600007ada000023efffffdc1100007adaffff8526ffffdc11;
    assign coff[1955] = 256'hffff8fb900003d76ffffc28affff8fb900007047ffffc28a00003d7600007047;
    assign coff[1956] = 256'h00006221ffffadd10000522f00006221ffff9ddf0000522fffffadd1ffff9ddf;
    assign coff[1957] = 256'hffff807ffffff4b900000b47ffff807f00007f8100000b47fffff4b900007f81;
    assign coff[1958] = 256'hffffd9a0ffff85e300007a1dffffd9a00000266000007a1dffff85e300002660;
    assign coff[1959] = 256'hffffc4ca0000717bffff8e85ffffc4ca00003b36ffff8e850000717b00003b36;
    assign coff[1960] = 256'h000075c3ffffcdd700003229000075c3ffff8a3d00003229ffffcdd7ffff8a3d;
    assign coff[1961] = 256'hffff8943ffffd03300002fcdffff8943000076bd00002fcdffffd033000076bd;
    assign coff[1962] = 256'hfffffeb9ffff800200007ffefffffeb90000014700007ffeffff800200000147;
    assign coff[1963] = 256'hffffa66600005b68ffffa498ffffa6660000599affffa49800005b680000599a;
    assign coff[1964] = 256'h0000460cffff94de00006b220000460cffffb9f400006b22ffff94deffffb9f4;
    assign coff[1965] = 256'hffff82b700001a39ffffe5c7ffff82b700007d49ffffe5c700001a3900007d49;
    assign coff[1966] = 256'hffffb7d4ffff9649000069b7ffffb7d40000482c000069b7ffff96490000482c;
    assign coff[1967] = 256'hffffe84800007dc9ffff8237ffffe848000017b8ffff823700007dc9000017b8;
    assign coff[1968] = 256'h00007bd9ffffdfa90000205700007bd9ffff842700002057ffffdfa9ffff8427;
    assign coff[1969] = 256'hffff918fffffbf4b000040b5ffff918f00006e71000040b5ffffbf4b00006e71;
    assign coff[1970] = 256'h00001185ffff813400007ecc00001185ffffee7b00007eccffff8134ffffee7b;
    assign coff[1971] = 256'hffff99f400004d45ffffb2bbffff99f40000660cffffb2bb00004d450000660c;
    assign coff[1972] = 256'h00005502ffffa04e00005fb200005502ffffaafe00005fb2ffffa04effffaafe;
    assign coff[1973] = 256'hffff80390000078efffff872ffff803900007fc7fffff8720000078e00007fc7;
    assign coff[1974] = 256'hffffc81fffff8cd700007329ffffc81f000037e100007329ffff8cd7000037e1;
    assign coff[1975] = 256'hffffd615000078f1ffff870fffffd615000029ebffff870f000078f1000029eb;
    assign coff[1976] = 256'h00006d21ffffbd1a000042e600006d21ffff92df000042e6ffffbd1affff92df;
    assign coff[1977] = 256'hffff8388ffffe22300001dddffff838800007c7800001dddffffe22300007c78;
    assign coff[1978] = 256'hffffebf5ffff819400007e6cffffebf50000140b00007e6cffff81940000140b;
    assign coff[1979] = 256'hffffb4c800006791ffff986fffffb4c800004b38ffff986f0000679100004b38;
    assign coff[1980] = 256'h00003592ffff8bc00000744000003592ffffca6e00007440ffff8bc0ffffca6e;
    assign coff[1981] = 256'hffff87eb00002c52ffffd3aeffff87eb00007815ffffd3ae00002c5200007815;
    assign coff[1982] = 256'hffffa919ffffa20500005dfbffffa919000056e700005dfbffffa205000056e7;
    assign coff[1983] = 256'hfffffaff00007fe7ffff8019fffffaff00000501ffff801900007fe700000501;
    assign coff[1984] = 256'h00007fadfffff6e10000091f00007fadffff80530000091ffffff6e1ffff8053;
    assign coff[1985] = 256'hffff9f45ffffac2c000053d4ffff9f45000060bb000053d4ffffac2c000060bb;
    assign coff[1986] = 256'h0000286effff868e000079720000286effffd79200007972ffff868effffd792;
    assign coff[1987] = 256'hffff8d8900003949ffffc6b7ffff8d8900007277ffffc6b70000394900007277;
    assign coff[1988] = 256'h00006517ffffb17c00004e8400006517ffff9ae900004e84ffffb17cffff9ae9;
    assign coff[1989] = 256'hffff8100fffff00a00000ff6ffff810000007f0000000ff6fffff00a00007f00;
    assign coff[1990] = 256'hffffde25ffff848f00007b71ffffde25000021db00007b71ffff848f000021db;
    assign coff[1991] = 256'hffffc0a700006f3affff90c6ffffc0a700003f59ffff90c600006f3a00003f59;
    assign coff[1992] = 256'h00007787ffffd23500002dcb00007787ffff887900002dcbffffd235ffff8879;
    assign coff[1993] = 256'hffff8b1affffcbdc00003424ffff8b1a000074e600003424ffffcbdc000074e6;
    assign coff[1994] = 256'h00000370ffff800c00007ff400000370fffffc9000007ff4ffff800cfffffc90;
    assign coff[1995] = 256'hffffa3180000580cffffa7f4ffffa31800005ce8ffffa7f40000580c00005ce8;
    assign coff[1996] = 256'h000049f2ffff97850000687b000049f2ffffb60e0000687bffff9785ffffb60e;
    assign coff[1997] = 256'hffff81d600001598ffffea68ffff81d600007e2affffea680000159800007e2a;
    assign coff[1998] = 256'hffffbbc5ffff93b400006c4cffffbbc50000443b00006c4cffff93b40000443b;
    assign coff[1999] = 256'hffffe3ab00007cd3ffff832dffffe3ab00001c55ffff832d00007cd300001c55;
    assign coff[2000] = 256'h00007cf4ffffe43e00001bc200007cf4ffff830c00001bc2ffffe43effff830c;
    assign coff[2001] = 256'hffff9404ffffbb46000044baffff940400006bfc000044baffffbb4600006bfc;
    assign coff[2002] = 256'h0000162cffff81ef00007e110000162cffffe9d400007e11ffff81efffffe9d4;
    assign coff[2003] = 256'hffff972e00004976ffffb68affff972e000068d2ffffb68a00004976000068d2;
    assign coff[2004] = 256'h00005879ffffa38000005c8000005879ffffa78700005c80ffffa380ffffa787;
    assign coff[2005] = 256'hffff8008000002d9fffffd27ffff800800007ff8fffffd27000002d900007ff8;
    assign coff[2006] = 256'hffffcc66ffff8add00007523ffffcc660000339a00007523ffff8add0000339a;
    assign coff[2007] = 256'hffffd1a900007751ffff88afffffd1a900002e57ffff88af0000775100002e57;
    assign coff[2008] = 256'h00006f84ffffc12a00003ed600006f84ffff907c00003ed6ffffc12affff907c;
    assign coff[2009] = 256'hffff84b7ffffdd940000226cffff84b700007b490000226cffffdd9400007b49;
    assign coff[2010] = 256'hfffff0a0ffff80ed00007f13fffff0a000000f6000007f13ffff80ed00000f60;
    assign coff[2011] = 256'hffffb105000064baffff9b46ffffb10500004efbffff9b46000064ba00004efb;
    assign coff[2012] = 256'h000039d0ffff8dcd00007233000039d0ffffc63000007233ffff8dcdffffc630;
    assign coff[2013] = 256'hffff865e000027dfffffd821ffff865e000079a2ffffd821000027df000079a2;
    assign coff[2014] = 256'hffffac9effff9ee30000611dffffac9e000053620000611dffff9ee300005362;
    assign coff[2015] = 256'hfffff64a00007fa2ffff805efffff64a000009b6ffff805e00007fa2000009b6;
    assign coff[2016] = 256'h00007ea8ffffed830000127d00007ea8ffff81580000127dffffed83ffff8158;
    assign coff[2017] = 256'hffff995dffffb38400004c7cffff995d000066a300004c7cffffb384000066a3;
    assign coff[2018] = 256'h00001f63ffff83e800007c1800001f63ffffe09d00007c18ffff83e8ffffe09d;
    assign coff[2019] = 256'hffff920f0000418dffffbe73ffff920f00006df1ffffbe730000418d00006df1;
    assign coff[2020] = 256'h00005f0affffaa42000055be00005f0affffa0f6000055beffffaa42ffffa0f6;
    assign coff[2021] = 256'hffff802bfffff96d00000693ffff802b00007fd500000693fffff96d00007fd5;
    assign coff[2022] = 256'hffffd528ffff87620000789effffd52800002ad80000789effff876200002ad8;
    assign coff[2023] = 256'hffffc90200007396ffff8c6affffc902000036feffff8c6a00007396000036fe;
    assign coff[2024] = 256'h000073d6ffffc98a00003676000073d6ffff8c2a00003676ffffc98affff8c2a;
    assign coff[2025] = 256'hffff8795ffffd49a00002b66ffff87950000786b00002b66ffffd49a0000786b;
    assign coff[2026] = 256'hfffffa03ffff802400007fdcfffffa03000005fd00007fdcffff8024000005fd;
    assign coff[2027] = 256'hffffa9d300005ea5ffffa15bffffa9d30000562dffffa15b00005ea50000562d;
    assign coff[2028] = 256'h0000420fffff925d00006da30000420fffffbdf100006da3ffff925dffffbdf1;
    assign coff[2029] = 256'hffff83c400001ed1ffffe12fffff83c400007c3cffffe12f00001ed100007c3c;
    assign coff[2030] = 256'hffffb3fdffff9904000066fcffffb3fd00004c03000066fcffff990400004c03;
    assign coff[2031] = 256'hffffeced00007e92ffff816effffeced00001313ffff816e00007e9200001313;
    assign coff[2032] = 256'h00007a93ffffdb20000024e000007a93ffff856d000024e0ffffdb20ffff856d;
    assign coff[2033] = 256'hffff8f41ffffc36700003c99ffff8f41000070bf00003c99ffffc367000070bf;
    assign coff[2034] = 256'h00000cd7ffff80a500007f5b00000cd7fffff32900007f5bffff80a5fffff329;
    assign coff[2035] = 256'hffff9cde000050f9ffffaf07ffff9cde00006322ffffaf07000050f900006322;
    assign coff[2036] = 256'h0000516effff9d3e000062c20000516effffae92000062c2ffff9d3effffae92;
    assign coff[2037] = 256'hffff809600000c41fffff3bfffff809600007f6afffff3bf00000c4100007f6a;
    assign coff[2038] = 256'hffffc3ecffff8efa00007106ffffc3ec00003c1400007106ffff8efa00003c14;
    assign coff[2039] = 256'hffffda9000007a67ffff8599ffffda9000002570ffff859900007a6700002570;
    assign coff[2040] = 256'h00006a97ffffb922000046de00006a97ffff9569000046deffffb922ffff9569;
    assign coff[2041] = 256'hffff8284ffffe6bd00001943ffff828400007d7c00001943ffffe6bd00007d7c;
    assign coff[2042] = 256'hffffe751ffff826700007d99ffffe751000018af00007d99ffff8267000018af;
    assign coff[2043] = 256'hffffb8a400006a44ffff95bcffffb8a40000475cffff95bc00006a440000475c;
    assign coff[2044] = 256'h00003141ffff89db0000762500003141ffffcebf00007625ffff89dbffffcebf;
    assign coff[2045] = 256'hffff89a2000030b6ffffcf4affff89a20000765effffcf4a000030b60000765e;
    assign coff[2046] = 256'hffffa5b3ffffa54800005ab8ffffa5b300005a4d00005ab8ffffa54800005a4d;
    assign coff[2047] = 256'hffffffb500007fffffff8001ffffffb50000004bffff800100007fff0000004b;

    always_ff @(posedge clk, negedge rst_n) begin
        if(~rst_n) begin
            data_o <= 'b0;
        end else if (valid == 1) begin
            data_o <= coff[addr_i];
        end else begin
            data_o <= 'b0;
        end
    end


endmodule