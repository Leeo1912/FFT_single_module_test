`timescale 1ns/1ps
module rom_1
(
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic                     valid,
    input  logic [10:0]              addr_i,
    output logic [255:0]             data_o
);

    logic [255:0] coff[2047:0];

    assign coff[0   ] = 256'h00007fff0000000000000000ffff8001ffff8001000000000000000000007fff;
    assign coff[1   ] = 256'h00005a82ffffa57effffa57effffa57effffa57e00005a8200005a8200005a82;
    assign coff[2   ] = 256'h00007642ffffcf04ffffcf04ffff89beffff89be000030fc000030fc00007642;
    assign coff[3   ] = 256'h000030fcffff89beffff89beffffcf04ffffcf040000764200007642000030fc;
    assign coff[4   ] = 256'h00007d8affffe707ffffe707ffff8276ffff8276000018f9000018f900007d8a;
    assign coff[5   ] = 256'h0000471dffff9592ffff9592ffffb8e3ffffb8e300006a6e00006a6e0000471d;
    assign coff[6   ] = 256'h00006a6effffb8e3ffffb8e3ffff9592ffff95920000471d0000471d00006a6e;
    assign coff[7   ] = 256'h000018f9ffff8276ffff8276ffffe707ffffe70700007d8a00007d8a000018f9;
    assign coff[8   ] = 256'h00007f62fffff374fffff374ffff809effff809e00000c8c00000c8c00007f62;
    assign coff[9   ] = 256'h00005134ffff9d0effff9d0effffaeccffffaecc000062f2000062f200005134;
    assign coff[10  ] = 256'h000070e3ffffc3a9ffffc3a9ffff8f1dffff8f1d00003c5700003c57000070e3;
    assign coff[11  ] = 256'h00002528ffff8583ffff8583ffffdad8ffffdad800007a7d00007a7d00002528;
    assign coff[12  ] = 256'h00007a7dffffdad8ffffdad8ffff8583ffff8583000025280000252800007a7d;
    assign coff[13  ] = 256'h00003c57ffff8f1dffff8f1dffffc3a9ffffc3a9000070e3000070e300003c57;
    assign coff[14  ] = 256'h000062f2ffffaeccffffaeccffff9d0effff9d0e0000513400005134000062f2;
    assign coff[15  ] = 256'h00000c8cffff809effff809efffff374fffff37400007f6200007f6200000c8c;
    assign coff[16  ] = 256'h00007fd9fffff9b8fffff9b8ffff8027ffff8027000006480000064800007fd9;
    assign coff[17  ] = 256'h000055f6ffffa129ffffa129ffffaa0affffaa0a00005ed700005ed7000055f6;
    assign coff[18  ] = 256'h000073b6ffffc946ffffc946ffff8c4affff8c4a000036ba000036ba000073b6;
    assign coff[19  ] = 256'h00002b1fffff877bffff877bffffd4e1ffffd4e1000078850000788500002b1f;
    assign coff[20  ] = 256'h00007c2affffe0e6ffffe0e6ffff83d6ffff83d600001f1a00001f1a00007c2a;
    assign coff[21  ] = 256'h000041ceffff9236ffff9236ffffbe32ffffbe3200006dca00006dca000041ce;
    assign coff[22  ] = 256'h000066d0ffffb3c0ffffb3c0ffff9930ffff993000004c4000004c40000066d0;
    assign coff[23  ] = 256'h000012c8ffff8163ffff8163ffffed38ffffed3800007e9d00007e9d000012c8;
    assign coff[24  ] = 256'h00007e9dffffed38ffffed38ffff8163ffff8163000012c8000012c800007e9d;
    assign coff[25  ] = 256'h00004c40ffff9930ffff9930ffffb3c0ffffb3c0000066d0000066d000004c40;
    assign coff[26  ] = 256'h00006dcaffffbe32ffffbe32ffff9236ffff9236000041ce000041ce00006dca;
    assign coff[27  ] = 256'h00001f1affff83d6ffff83d6ffffe0e6ffffe0e600007c2a00007c2a00001f1a;
    assign coff[28  ] = 256'h00007885ffffd4e1ffffd4e1ffff877bffff877b00002b1f00002b1f00007885;
    assign coff[29  ] = 256'h000036baffff8c4affff8c4affffc946ffffc946000073b6000073b6000036ba;
    assign coff[30  ] = 256'h00005ed7ffffaa0affffaa0affffa129ffffa129000055f6000055f600005ed7;
    assign coff[31  ] = 256'h00000648ffff8027ffff8027fffff9b8fffff9b800007fd900007fd900000648;
    assign coff[32  ] = 256'h00007ff6fffffcdcfffffcdcffff800affff800a000003240000032400007ff6;
    assign coff[33  ] = 256'h00005843ffffa34cffffa34cffffa7bdffffa7bd00005cb400005cb400005843;
    assign coff[34  ] = 256'h00007505ffffcc21ffffcc21ffff8afbffff8afb000033df000033df00007505;
    assign coff[35  ] = 256'h00002e11ffff8894ffff8894ffffd1efffffd1ef0000776c0000776c00002e11;
    assign coff[36  ] = 256'h00007ce4ffffe3f4ffffe3f4ffff831cffff831c00001c0c00001c0c00007ce4;
    assign coff[37  ] = 256'h0000447bffff93dcffff93dcffffbb85ffffbb8500006c2400006c240000447b;
    assign coff[38  ] = 256'h000068a7ffffb64cffffb64cffff9759ffff9759000049b4000049b4000068a7;
    assign coff[39  ] = 256'h000015e2ffff81e2ffff81e2ffffea1effffea1e00007e1e00007e1e000015e2;
    assign coff[40  ] = 256'h00007f0afffff055fffff055ffff80f6ffff80f600000fab00000fab00007f0a;
    assign coff[41  ] = 256'h00004ec0ffff9b17ffff9b17ffffb140ffffb140000064e9000064e900004ec0;
    assign coff[42  ] = 256'h00006f5fffffc0e9ffffc0e9ffff90a1ffff90a100003f1700003f1700006f5f;
    assign coff[43  ] = 256'h00002224ffff84a3ffff84a3ffffdddcffffdddc00007b5d00007b5d00002224;
    assign coff[44  ] = 256'h0000798affffd7d9ffffd7d9ffff8676ffff867600002827000028270000798a;
    assign coff[45  ] = 256'h0000398dffff8dabffff8dabffffc673ffffc67300007255000072550000398d;
    assign coff[46  ] = 256'h000060ecffffac65ffffac65ffff9f14ffff9f140000539b0000539b000060ec;
    assign coff[47  ] = 256'h0000096bffff8059ffff8059fffff695fffff69500007fa700007fa70000096b;
    assign coff[48  ] = 256'h00007fa7fffff695fffff695ffff8059ffff80590000096b0000096b00007fa7;
    assign coff[49  ] = 256'h0000539bffff9f14ffff9f14ffffac65ffffac65000060ec000060ec0000539b;
    assign coff[50  ] = 256'h00007255ffffc673ffffc673ffff8dabffff8dab0000398d0000398d00007255;
    assign coff[51  ] = 256'h00002827ffff8676ffff8676ffffd7d9ffffd7d90000798a0000798a00002827;
    assign coff[52  ] = 256'h00007b5dffffdddcffffdddcffff84a3ffff84a3000022240000222400007b5d;
    assign coff[53  ] = 256'h00003f17ffff90a1ffff90a1ffffc0e9ffffc0e900006f5f00006f5f00003f17;
    assign coff[54  ] = 256'h000064e9ffffb140ffffb140ffff9b17ffff9b1700004ec000004ec0000064e9;
    assign coff[55  ] = 256'h00000fabffff80f6ffff80f6fffff055fffff05500007f0a00007f0a00000fab;
    assign coff[56  ] = 256'h00007e1effffea1effffea1effff81e2ffff81e2000015e2000015e200007e1e;
    assign coff[57  ] = 256'h000049b4ffff9759ffff9759ffffb64cffffb64c000068a7000068a7000049b4;
    assign coff[58  ] = 256'h00006c24ffffbb85ffffbb85ffff93dcffff93dc0000447b0000447b00006c24;
    assign coff[59  ] = 256'h00001c0cffff831cffff831cffffe3f4ffffe3f400007ce400007ce400001c0c;
    assign coff[60  ] = 256'h0000776cffffd1efffffd1efffff8894ffff889400002e1100002e110000776c;
    assign coff[61  ] = 256'h000033dfffff8afbffff8afbffffcc21ffffcc210000750500007505000033df;
    assign coff[62  ] = 256'h00005cb4ffffa7bdffffa7bdffffa34cffffa34c000058430000584300005cb4;
    assign coff[63  ] = 256'h00000324ffff800affff800afffffcdcfffffcdc00007ff600007ff600000324;
    assign coff[64  ] = 256'h00007ffefffffe6efffffe6effff8002ffff8002000001920000019200007ffe;
    assign coff[65  ] = 256'h00005964ffffa463ffffa463ffffa69cffffa69c00005b9d00005b9d00005964;
    assign coff[66  ] = 256'h000075a6ffffcd92ffffcd92ffff8a5affff8a5a0000326e0000326e000075a6;
    assign coff[67  ] = 256'h00002f87ffff8927ffff8927ffffd079ffffd079000076d9000076d900002f87;
    assign coff[68  ] = 256'h00007d3affffe57dffffe57dffff82c6ffff82c600001a8300001a8300007d3a;
    assign coff[69  ] = 256'h000045cdffff94b5ffff94b5ffffba33ffffba3300006b4b00006b4b000045cd;
    assign coff[70  ] = 256'h0000698cffffb796ffffb796ffff9674ffff96740000486a0000486a0000698c;
    assign coff[71  ] = 256'h0000176effff822affff822affffe892ffffe89200007dd600007dd60000176e;
    assign coff[72  ] = 256'h00007f38fffff1e4fffff1e4ffff80c8ffff80c800000e1c00000e1c00007f38;
    assign coff[73  ] = 256'h00004ffbffff9c11ffff9c11ffffb005ffffb005000063ef000063ef00004ffb;
    assign coff[74  ] = 256'h00007023ffffc248ffffc248ffff8fddffff8fdd00003db800003db800007023;
    assign coff[75  ] = 256'h000023a7ffff8511ffff8511ffffdc59ffffdc5900007aef00007aef000023a7;
    assign coff[76  ] = 256'h00007a06ffffd958ffffd958ffff85faffff85fa000026a8000026a800007a06;
    assign coff[77  ] = 256'h00003af3ffff8e62ffff8e62ffffc50dffffc50d0000719e0000719e00003af3;
    assign coff[78  ] = 256'h000061f1ffffad97ffffad97ffff9e0fffff9e0f0000526900005269000061f1;
    assign coff[79  ] = 256'h00000afbffff8079ffff8079fffff505fffff50500007f8700007f8700000afb;
    assign coff[80  ] = 256'h00007fc2fffff827fffff827ffff803effff803e000007d9000007d900007fc2;
    assign coff[81  ] = 256'h000054caffffa01cffffa01cffffab36ffffab3600005fe400005fe4000054ca;
    assign coff[82  ] = 256'h00007308ffffc7dbffffc7dbffff8cf8ffff8cf8000038250000382500007308;
    assign coff[83  ] = 256'h000029a4ffff86f6ffff86f6ffffd65cffffd65c0000790a0000790a000029a4;
    assign coff[84  ] = 256'h00007bc6ffffdf61ffffdf61ffff843affff843a0000209f0000209f00007bc6;
    assign coff[85  ] = 256'h00004074ffff9169ffff9169ffffbf8cffffbf8c00006e9700006e9700004074;
    assign coff[86  ] = 256'h000065deffffb27fffffb27fffff9a22ffff9a2200004d8100004d81000065de;
    assign coff[87  ] = 256'h0000113affff812affff812affffeec6ffffeec600007ed600007ed60000113a;
    assign coff[88  ] = 256'h00007e60ffffebabffffebabffff81a0ffff81a0000014550000145500007e60;
    assign coff[89  ] = 256'h00004afbffff9843ffff9843ffffb505ffffb505000067bd000067bd00004afb;
    assign coff[90  ] = 256'h00006cf9ffffbcdaffffbcdaffff9307ffff9307000043260000432600006cf9;
    assign coff[91  ] = 256'h00001d93ffff8377ffff8377ffffe26dffffe26d00007c8900007c8900001d93;
    assign coff[92  ] = 256'h000077fbffffd367ffffd367ffff8805ffff880500002c9900002c99000077fb;
    assign coff[93  ] = 256'h0000354effff8ba0ffff8ba0ffffcab2ffffcab200007460000074600000354e;
    assign coff[94  ] = 256'h00005dc8ffffa8e2ffffa8e2ffffa238ffffa2380000571e0000571e00005dc8;
    assign coff[95  ] = 256'h000004b6ffff8016ffff8016fffffb4afffffb4a00007fea00007fea000004b6;
    assign coff[96  ] = 256'h00007feafffffb4afffffb4affff8016ffff8016000004b6000004b600007fea;
    assign coff[97  ] = 256'h0000571effffa238ffffa238ffffa8e2ffffa8e200005dc800005dc80000571e;
    assign coff[98  ] = 256'h00007460ffffcab2ffffcab2ffff8ba0ffff8ba00000354e0000354e00007460;
    assign coff[99  ] = 256'h00002c99ffff8805ffff8805ffffd367ffffd367000077fb000077fb00002c99;
    assign coff[100 ] = 256'h00007c89ffffe26dffffe26dffff8377ffff837700001d9300001d9300007c89;
    assign coff[101 ] = 256'h00004326ffff9307ffff9307ffffbcdaffffbcda00006cf900006cf900004326;
    assign coff[102 ] = 256'h000067bdffffb505ffffb505ffff9843ffff984300004afb00004afb000067bd;
    assign coff[103 ] = 256'h00001455ffff81a0ffff81a0ffffebabffffebab00007e6000007e6000001455;
    assign coff[104 ] = 256'h00007ed6ffffeec6ffffeec6ffff812affff812a0000113a0000113a00007ed6;
    assign coff[105 ] = 256'h00004d81ffff9a22ffff9a22ffffb27fffffb27f000065de000065de00004d81;
    assign coff[106 ] = 256'h00006e97ffffbf8cffffbf8cffff9169ffff9169000040740000407400006e97;
    assign coff[107 ] = 256'h0000209fffff843affff843affffdf61ffffdf6100007bc600007bc60000209f;
    assign coff[108 ] = 256'h0000790affffd65cffffd65cffff86f6ffff86f6000029a4000029a40000790a;
    assign coff[109 ] = 256'h00003825ffff8cf8ffff8cf8ffffc7dbffffc7db000073080000730800003825;
    assign coff[110 ] = 256'h00005fe4ffffab36ffffab36ffffa01cffffa01c000054ca000054ca00005fe4;
    assign coff[111 ] = 256'h000007d9ffff803effff803efffff827fffff82700007fc200007fc2000007d9;
    assign coff[112 ] = 256'h00007f87fffff505fffff505ffff8079ffff807900000afb00000afb00007f87;
    assign coff[113 ] = 256'h00005269ffff9e0fffff9e0fffffad97ffffad97000061f1000061f100005269;
    assign coff[114 ] = 256'h0000719effffc50dffffc50dffff8e62ffff8e6200003af300003af30000719e;
    assign coff[115 ] = 256'h000026a8ffff85faffff85faffffd958ffffd95800007a0600007a06000026a8;
    assign coff[116 ] = 256'h00007aefffffdc59ffffdc59ffff8511ffff8511000023a7000023a700007aef;
    assign coff[117 ] = 256'h00003db8ffff8fddffff8fddffffc248ffffc248000070230000702300003db8;
    assign coff[118 ] = 256'h000063efffffb005ffffb005ffff9c11ffff9c1100004ffb00004ffb000063ef;
    assign coff[119 ] = 256'h00000e1cffff80c8ffff80c8fffff1e4fffff1e400007f3800007f3800000e1c;
    assign coff[120 ] = 256'h00007dd6ffffe892ffffe892ffff822affff822a0000176e0000176e00007dd6;
    assign coff[121 ] = 256'h0000486affff9674ffff9674ffffb796ffffb7960000698c0000698c0000486a;
    assign coff[122 ] = 256'h00006b4bffffba33ffffba33ffff94b5ffff94b5000045cd000045cd00006b4b;
    assign coff[123 ] = 256'h00001a83ffff82c6ffff82c6ffffe57dffffe57d00007d3a00007d3a00001a83;
    assign coff[124 ] = 256'h000076d9ffffd079ffffd079ffff8927ffff892700002f8700002f87000076d9;
    assign coff[125 ] = 256'h0000326effff8a5affff8a5affffcd92ffffcd92000075a6000075a60000326e;
    assign coff[126 ] = 256'h00005b9dffffa69cffffa69cffffa463ffffa463000059640000596400005b9d;
    assign coff[127 ] = 256'h00000192ffff8002ffff8002fffffe6efffffe6e00007ffe00007ffe00000192;
    assign coff[128 ] = 256'h00007fffffffff37ffffff37ffff8001ffff8001000000c9000000c900007fff;
    assign coff[129 ] = 256'h000059f4ffffa4f0ffffa4f0ffffa60cffffa60c00005b1000005b10000059f4;
    assign coff[130 ] = 256'h000075f4ffffce4bffffce4bffff8a0cffff8a0c000031b5000031b5000075f4;
    assign coff[131 ] = 256'h00003042ffff8972ffff8972ffffcfbeffffcfbe0000768e0000768e00003042;
    assign coff[132 ] = 256'h00007d63ffffe642ffffe642ffff829dffff829d000019be000019be00007d63;
    assign coff[133 ] = 256'h00004675ffff9523ffff9523ffffb98bffffb98b00006add00006add00004675;
    assign coff[134 ] = 256'h000069fdffffb83cffffb83cffff9603ffff9603000047c4000047c4000069fd;
    assign coff[135 ] = 256'h00001833ffff824fffff824fffffe7cdffffe7cd00007db100007db100001833;
    assign coff[136 ] = 256'h00007f4efffff2acfffff2acffff80b2ffff80b200000d5400000d5400007f4e;
    assign coff[137 ] = 256'h00005098ffff9c8fffff9c8fffffaf68ffffaf68000063710000637100005098;
    assign coff[138 ] = 256'h00007083ffffc2f8ffffc2f8ffff8f7dffff8f7d00003d0800003d0800007083;
    assign coff[139 ] = 256'h00002467ffff8549ffff8549ffffdb99ffffdb9900007ab700007ab700002467;
    assign coff[140 ] = 256'h00007a42ffffda18ffffda18ffff85beffff85be000025e8000025e800007a42;
    assign coff[141 ] = 256'h00003ba5ffff8ebfffff8ebfffffc45bffffc45b000071410000714100003ba5;
    assign coff[142 ] = 256'h00006272ffffae31ffffae31ffff9d8effff9d8e000051cf000051cf00006272;
    assign coff[143 ] = 256'h00000bc4ffff808bffff808bfffff43cfffff43c00007f7500007f7500000bc4;
    assign coff[144 ] = 256'h00007fcefffff8effffff8efffff8032ffff8032000007110000071100007fce;
    assign coff[145 ] = 256'h00005560ffffa0a2ffffa0a2ffffaaa0ffffaaa000005f5e00005f5e00005560;
    assign coff[146 ] = 256'h0000735fffffc890ffffc890ffff8ca1ffff8ca100003770000037700000735f;
    assign coff[147 ] = 256'h00002a62ffff8738ffff8738ffffd59effffd59e000078c8000078c800002a62;
    assign coff[148 ] = 256'h00007bf9ffffe023ffffe023ffff8407ffff840700001fdd00001fdd00007bf9;
    assign coff[149 ] = 256'h00004121ffff91cfffff91cfffffbedfffffbedf00006e3100006e3100004121;
    assign coff[150 ] = 256'h00006657ffffb31fffffb31fffff99a9ffff99a900004ce100004ce100006657;
    assign coff[151 ] = 256'h00001201ffff8146ffff8146ffffedffffffedff00007eba00007eba00001201;
    assign coff[152 ] = 256'h00007e7fffffec71ffffec71ffff8181ffff81810000138f0000138f00007e7f;
    assign coff[153 ] = 256'h00004b9effff98b9ffff98b9ffffb462ffffb462000067470000674700004b9e;
    assign coff[154 ] = 256'h00006d62ffffbd86ffffbd86ffff929effff929e0000427a0000427a00006d62;
    assign coff[155 ] = 256'h00001e57ffff83a6ffff83a6ffffe1a9ffffe1a900007c5a00007c5a00001e57;
    assign coff[156 ] = 256'h00007840ffffd424ffffd424ffff87c0ffff87c000002bdc00002bdc00007840;
    assign coff[157 ] = 256'h00003604ffff8bf5ffff8bf5ffffc9fcffffc9fc0000740b0000740b00003604;
    assign coff[158 ] = 256'h00005e50ffffa976ffffa976ffffa1b0ffffa1b00000568a0000568a00005e50;
    assign coff[159 ] = 256'h0000057fffff801effff801efffffa81fffffa8100007fe200007fe20000057f;
    assign coff[160 ] = 256'h00007ff1fffffc13fffffc13ffff800fffff800f000003ed000003ed00007ff1;
    assign coff[161 ] = 256'h000057b1ffffa2c2ffffa2c2ffffa84fffffa84f00005d3e00005d3e000057b1;
    assign coff[162 ] = 256'h000074b3ffffcb69ffffcb69ffff8b4dffff8b4d0000349700003497000074b3;
    assign coff[163 ] = 256'h00002d55ffff884cffff884cffffd2abffffd2ab000077b4000077b400002d55;
    assign coff[164 ] = 256'h00007cb7ffffe330ffffe330ffff8349ffff834900001cd000001cd000007cb7;
    assign coff[165 ] = 256'h000043d1ffff9371ffff9371ffffbc2fffffbc2f00006c8f00006c8f000043d1;
    assign coff[166 ] = 256'h00006832ffffb5a8ffffb5a8ffff97ceffff97ce00004a5800004a5800006832;
    assign coff[167 ] = 256'h0000151cffff81c1ffff81c1ffffeae4ffffeae400007e3f00007e3f0000151c;
    assign coff[168 ] = 256'h00007ef0ffffef8dffffef8dffff8110ffff8110000010730000107300007ef0;
    assign coff[169 ] = 256'h00004e21ffff9a9cffff9a9cffffb1dfffffb1df000065640000656400004e21;
    assign coff[170 ] = 256'h00006efbffffc03affffc03affff9105ffff910500003fc600003fc600006efb;
    assign coff[171 ] = 256'h00002162ffff846effff846effffde9effffde9e00007b9200007b9200002162;
    assign coff[172 ] = 256'h0000794affffd71bffffd71bffff86b6ffff86b6000028e5000028e50000794a;
    assign coff[173 ] = 256'h000038d9ffff8d51ffff8d51ffffc727ffffc727000072af000072af000038d9;
    assign coff[174 ] = 256'h00006068ffffabcdffffabcdffff9f98ffff9f98000054330000543300006068;
    assign coff[175 ] = 256'h000008a2ffff804bffff804bfffff75efffff75e00007fb500007fb5000008a2;
    assign coff[176 ] = 256'h00007f98fffff5cdfffff5cdffff8068ffff806800000a3300000a3300007f98;
    assign coff[177 ] = 256'h00005303ffff9e91ffff9e91ffffacfdffffacfd0000616f0000616f00005303;
    assign coff[178 ] = 256'h000071faffffc5c0ffffc5c0ffff8e06ffff8e0600003a4000003a40000071fa;
    assign coff[179 ] = 256'h00002768ffff8637ffff8637ffffd898ffffd898000079c9000079c900002768;
    assign coff[180 ] = 256'h00007b27ffffdd1bffffdd1bffff84d9ffff84d9000022e5000022e500007b27;
    assign coff[181 ] = 256'h00003e68ffff903effff903effffc198ffffc19800006fc200006fc200003e68;
    assign coff[182 ] = 256'h0000646cffffb0a2ffffb0a2ffff9b94ffff9b9400004f5e00004f5e0000646c;
    assign coff[183 ] = 256'h00000ee4ffff80deffff80defffff11cfffff11c00007f2200007f2200000ee4;
    assign coff[184 ] = 256'h00007dfbffffe958ffffe958ffff8205ffff8205000016a8000016a800007dfb;
    assign coff[185 ] = 256'h0000490fffff96e6ffff96e6ffffb6f1ffffb6f10000691a0000691a0000490f;
    assign coff[186 ] = 256'h00006bb8ffffbadcffffbadcffff9448ffff9448000045240000452400006bb8;
    assign coff[187 ] = 256'h00001b47ffff82f1ffff82f1ffffe4b9ffffe4b900007d0f00007d0f00001b47;
    assign coff[188 ] = 256'h00007723ffffd134ffffd134ffff88ddffff88dd00002ecc00002ecc00007723;
    assign coff[189 ] = 256'h00003327ffff8aaaffff8aaaffffccd9ffffccd9000075560000755600003327;
    assign coff[190 ] = 256'h00005c29ffffa72cffffa72cffffa3d7ffffa3d7000058d4000058d400005c29;
    assign coff[191 ] = 256'h0000025bffff8006ffff8006fffffda5fffffda500007ffa00007ffa0000025b;
    assign coff[192 ] = 256'h00007ffafffffda5fffffda5ffff8006ffff80060000025b0000025b00007ffa;
    assign coff[193 ] = 256'h000058d4ffffa3d7ffffa3d7ffffa72cffffa72c00005c2900005c29000058d4;
    assign coff[194 ] = 256'h00007556ffffccd9ffffccd9ffff8aaaffff8aaa000033270000332700007556;
    assign coff[195 ] = 256'h00002eccffff88ddffff88ddffffd134ffffd134000077230000772300002ecc;
    assign coff[196 ] = 256'h00007d0fffffe4b9ffffe4b9ffff82f1ffff82f100001b4700001b4700007d0f;
    assign coff[197 ] = 256'h00004524ffff9448ffff9448ffffbadcffffbadc00006bb800006bb800004524;
    assign coff[198 ] = 256'h0000691affffb6f1ffffb6f1ffff96e6ffff96e60000490f0000490f0000691a;
    assign coff[199 ] = 256'h000016a8ffff8205ffff8205ffffe958ffffe95800007dfb00007dfb000016a8;
    assign coff[200 ] = 256'h00007f22fffff11cfffff11cffff80deffff80de00000ee400000ee400007f22;
    assign coff[201 ] = 256'h00004f5effff9b94ffff9b94ffffb0a2ffffb0a20000646c0000646c00004f5e;
    assign coff[202 ] = 256'h00006fc2ffffc198ffffc198ffff903effff903e00003e6800003e6800006fc2;
    assign coff[203 ] = 256'h000022e5ffff84d9ffff84d9ffffdd1bffffdd1b00007b2700007b27000022e5;
    assign coff[204 ] = 256'h000079c9ffffd898ffffd898ffff8637ffff86370000276800002768000079c9;
    assign coff[205 ] = 256'h00003a40ffff8e06ffff8e06ffffc5c0ffffc5c0000071fa000071fa00003a40;
    assign coff[206 ] = 256'h0000616fffffacfdffffacfdffff9e91ffff9e9100005303000053030000616f;
    assign coff[207 ] = 256'h00000a33ffff8068ffff8068fffff5cdfffff5cd00007f9800007f9800000a33;
    assign coff[208 ] = 256'h00007fb5fffff75efffff75effff804bffff804b000008a2000008a200007fb5;
    assign coff[209 ] = 256'h00005433ffff9f98ffff9f98ffffabcdffffabcd000060680000606800005433;
    assign coff[210 ] = 256'h000072afffffc727ffffc727ffff8d51ffff8d51000038d9000038d9000072af;
    assign coff[211 ] = 256'h000028e5ffff86b6ffff86b6ffffd71bffffd71b0000794a0000794a000028e5;
    assign coff[212 ] = 256'h00007b92ffffde9effffde9effff846effff846e000021620000216200007b92;
    assign coff[213 ] = 256'h00003fc6ffff9105ffff9105ffffc03affffc03a00006efb00006efb00003fc6;
    assign coff[214 ] = 256'h00006564ffffb1dfffffb1dfffff9a9cffff9a9c00004e2100004e2100006564;
    assign coff[215 ] = 256'h00001073ffff8110ffff8110ffffef8dffffef8d00007ef000007ef000001073;
    assign coff[216 ] = 256'h00007e3fffffeae4ffffeae4ffff81c1ffff81c10000151c0000151c00007e3f;
    assign coff[217 ] = 256'h00004a58ffff97ceffff97ceffffb5a8ffffb5a8000068320000683200004a58;
    assign coff[218 ] = 256'h00006c8fffffbc2fffffbc2fffff9371ffff9371000043d1000043d100006c8f;
    assign coff[219 ] = 256'h00001cd0ffff8349ffff8349ffffe330ffffe33000007cb700007cb700001cd0;
    assign coff[220 ] = 256'h000077b4ffffd2abffffd2abffff884cffff884c00002d5500002d55000077b4;
    assign coff[221 ] = 256'h00003497ffff8b4dffff8b4dffffcb69ffffcb69000074b3000074b300003497;
    assign coff[222 ] = 256'h00005d3effffa84fffffa84fffffa2c2ffffa2c2000057b1000057b100005d3e;
    assign coff[223 ] = 256'h000003edffff800fffff800ffffffc13fffffc1300007ff100007ff1000003ed;
    assign coff[224 ] = 256'h00007fe2fffffa81fffffa81ffff801effff801e0000057f0000057f00007fe2;
    assign coff[225 ] = 256'h0000568affffa1b0ffffa1b0ffffa976ffffa97600005e5000005e500000568a;
    assign coff[226 ] = 256'h0000740bffffc9fcffffc9fcffff8bf5ffff8bf500003604000036040000740b;
    assign coff[227 ] = 256'h00002bdcffff87c0ffff87c0ffffd424ffffd424000078400000784000002bdc;
    assign coff[228 ] = 256'h00007c5affffe1a9ffffe1a9ffff83a6ffff83a600001e5700001e5700007c5a;
    assign coff[229 ] = 256'h0000427affff929effff929effffbd86ffffbd8600006d6200006d620000427a;
    assign coff[230 ] = 256'h00006747ffffb462ffffb462ffff98b9ffff98b900004b9e00004b9e00006747;
    assign coff[231 ] = 256'h0000138fffff8181ffff8181ffffec71ffffec7100007e7f00007e7f0000138f;
    assign coff[232 ] = 256'h00007ebaffffedffffffedffffff8146ffff8146000012010000120100007eba;
    assign coff[233 ] = 256'h00004ce1ffff99a9ffff99a9ffffb31fffffb31f000066570000665700004ce1;
    assign coff[234 ] = 256'h00006e31ffffbedfffffbedfffff91cfffff91cf000041210000412100006e31;
    assign coff[235 ] = 256'h00001fddffff8407ffff8407ffffe023ffffe02300007bf900007bf900001fdd;
    assign coff[236 ] = 256'h000078c8ffffd59effffd59effff8738ffff873800002a6200002a62000078c8;
    assign coff[237 ] = 256'h00003770ffff8ca1ffff8ca1ffffc890ffffc8900000735f0000735f00003770;
    assign coff[238 ] = 256'h00005f5effffaaa0ffffaaa0ffffa0a2ffffa0a2000055600000556000005f5e;
    assign coff[239 ] = 256'h00000711ffff8032ffff8032fffff8effffff8ef00007fce00007fce00000711;
    assign coff[240 ] = 256'h00007f75fffff43cfffff43cffff808bffff808b00000bc400000bc400007f75;
    assign coff[241 ] = 256'h000051cfffff9d8effff9d8effffae31ffffae310000627200006272000051cf;
    assign coff[242 ] = 256'h00007141ffffc45bffffc45bffff8ebfffff8ebf00003ba500003ba500007141;
    assign coff[243 ] = 256'h000025e8ffff85beffff85beffffda18ffffda1800007a4200007a42000025e8;
    assign coff[244 ] = 256'h00007ab7ffffdb99ffffdb99ffff8549ffff8549000024670000246700007ab7;
    assign coff[245 ] = 256'h00003d08ffff8f7dffff8f7dffffc2f8ffffc2f8000070830000708300003d08;
    assign coff[246 ] = 256'h00006371ffffaf68ffffaf68ffff9c8fffff9c8f000050980000509800006371;
    assign coff[247 ] = 256'h00000d54ffff80b2ffff80b2fffff2acfffff2ac00007f4e00007f4e00000d54;
    assign coff[248 ] = 256'h00007db1ffffe7cdffffe7cdffff824fffff824f000018330000183300007db1;
    assign coff[249 ] = 256'h000047c4ffff9603ffff9603ffffb83cffffb83c000069fd000069fd000047c4;
    assign coff[250 ] = 256'h00006addffffb98bffffb98bffff9523ffff9523000046750000467500006add;
    assign coff[251 ] = 256'h000019beffff829dffff829dffffe642ffffe64200007d6300007d63000019be;
    assign coff[252 ] = 256'h0000768effffcfbeffffcfbeffff8972ffff897200003042000030420000768e;
    assign coff[253 ] = 256'h000031b5ffff8a0cffff8a0cffffce4bffffce4b000075f4000075f4000031b5;
    assign coff[254 ] = 256'h00005b10ffffa60cffffa60cffffa4f0ffffa4f0000059f4000059f400005b10;
    assign coff[255 ] = 256'h000000c9ffff8001ffff8001ffffff37ffffff3700007fff00007fff000000c9;
    assign coff[256 ] = 256'h00007fffffffff9bffffff9bffff8001ffff8001000000650000006500007fff;
    assign coff[257 ] = 256'h00005a3bffffa537ffffa537ffffa5c5ffffa5c500005ac900005ac900005a3b;
    assign coff[258 ] = 256'h0000761bffffcea7ffffcea7ffff89e5ffff89e500003159000031590000761b;
    assign coff[259 ] = 256'h0000309fffff8998ffff8998ffffcf61ffffcf6100007668000076680000309f;
    assign coff[260 ] = 256'h00007d77ffffe6a5ffffe6a5ffff8289ffff82890000195b0000195b00007d77;
    assign coff[261 ] = 256'h000046c9ffff955bffff955bffffb937ffffb93700006aa500006aa5000046c9;
    assign coff[262 ] = 256'h00006a36ffffb890ffffb890ffff95caffff95ca000047700000477000006a36;
    assign coff[263 ] = 256'h00001896ffff8262ffff8262ffffe76affffe76a00007d9e00007d9e00001896;
    assign coff[264 ] = 256'h00007f58fffff310fffff310ffff80a8ffff80a800000cf000000cf000007f58;
    assign coff[265 ] = 256'h000050e6ffff9cceffff9cceffffaf1affffaf1a0000633200006332000050e6;
    assign coff[266 ] = 256'h000070b3ffffc351ffffc351ffff8f4dffff8f4d00003caf00003caf000070b3;
    assign coff[267 ] = 256'h000024c8ffff8566ffff8566ffffdb38ffffdb3800007a9a00007a9a000024c8;
    assign coff[268 ] = 256'h00007a60ffffda78ffffda78ffff85a0ffff85a0000025880000258800007a60;
    assign coff[269 ] = 256'h00003bfeffff8eeeffff8eeeffffc402ffffc402000071120000711200003bfe;
    assign coff[270 ] = 256'h000062b2ffffae7fffffae7fffff9d4effff9d4e0000518100005181000062b2;
    assign coff[271 ] = 256'h00000c28ffff8094ffff8094fffff3d8fffff3d800007f6c00007f6c00000c28;
    assign coff[272 ] = 256'h00007fd3fffff954fffff954ffff802dffff802d000006ac000006ac00007fd3;
    assign coff[273 ] = 256'h000055abffffa0e5ffffa0e5ffffaa55ffffaa5500005f1b00005f1b000055ab;
    assign coff[274 ] = 256'h0000738bffffc8ebffffc8ebffff8c75ffff8c7500003715000037150000738b;
    assign coff[275 ] = 256'h00002ac1ffff875affff875affffd53fffffd53f000078a6000078a600002ac1;
    assign coff[276 ] = 256'h00007c11ffffe085ffffe085ffff83efffff83ef00001f7b00001f7b00007c11;
    assign coff[277 ] = 256'h00004178ffff9202ffff9202ffffbe88ffffbe8800006dfe00006dfe00004178;
    assign coff[278 ] = 256'h00006693ffffb36fffffb36fffff996dffff996d00004c9100004c9100006693;
    assign coff[279 ] = 256'h00001265ffff8154ffff8154ffffed9bffffed9b00007eac00007eac00001265;
    assign coff[280 ] = 256'h00007e8effffecd5ffffecd5ffff8172ffff81720000132b0000132b00007e8e;
    assign coff[281 ] = 256'h00004befffff98f5ffff98f5ffffb411ffffb4110000670b0000670b00004bef;
    assign coff[282 ] = 256'h00006d96ffffbddcffffbddcffff926affff926a000042240000422400006d96;
    assign coff[283 ] = 256'h00001eb8ffff83beffff83beffffe148ffffe14800007c4200007c4200001eb8;
    assign coff[284 ] = 256'h00007863ffffd482ffffd482ffff879dffff879d00002b7e00002b7e00007863;
    assign coff[285 ] = 256'h0000365fffff8c1fffff8c1fffffc9a1ffffc9a1000073e1000073e10000365f;
    assign coff[286 ] = 256'h00005e94ffffa9c0ffffa9c0ffffa16cffffa16c000056400000564000005e94;
    assign coff[287 ] = 256'h000005e3ffff8023ffff8023fffffa1dfffffa1d00007fdd00007fdd000005e3;
    assign coff[288 ] = 256'h00007ff4fffffc77fffffc77ffff800cffff800c000003890000038900007ff4;
    assign coff[289 ] = 256'h000057faffffa307ffffa307ffffa806ffffa80600005cf900005cf9000057fa;
    assign coff[290 ] = 256'h000074dcffffcbc5ffffcbc5ffff8b24ffff8b240000343b0000343b000074dc;
    assign coff[291 ] = 256'h00002db3ffff8870ffff8870ffffd24dffffd24d000077900000779000002db3;
    assign coff[292 ] = 256'h00007cceffffe392ffffe392ffff8332ffff833200001c6e00001c6e00007cce;
    assign coff[293 ] = 256'h00004426ffff93a6ffff93a6ffffbbdaffffbbda00006c5a00006c5a00004426;
    assign coff[294 ] = 256'h0000686dffffb5faffffb5faffff9793ffff979300004a0600004a060000686d;
    assign coff[295 ] = 256'h0000157fffff81d1ffff81d1ffffea81ffffea8100007e2f00007e2f0000157f;
    assign coff[296 ] = 256'h00007efdffffeff1ffffeff1ffff8103ffff81030000100f0000100f00007efd;
    assign coff[297 ] = 256'h00004e71ffff9adaffff9adaffffb18fffffb18f000065260000652600004e71;
    assign coff[298 ] = 256'h00006f2dffffc091ffffc091ffff90d3ffff90d300003f6f00003f6f00006f2d;
    assign coff[299 ] = 256'h000021c3ffff8488ffff8488ffffde3dffffde3d00007b7800007b78000021c3;
    assign coff[300 ] = 256'h0000796affffd77affffd77affff8696ffff869600002886000028860000796a;
    assign coff[301 ] = 256'h00003933ffff8d7effff8d7effffc6cdffffc6cd000072820000728200003933;
    assign coff[302 ] = 256'h000060aaffffac19ffffac19ffff9f56ffff9f56000053e7000053e7000060aa;
    assign coff[303 ] = 256'h00000906ffff8052ffff8052fffff6fafffff6fa00007fae00007fae00000906;
    assign coff[304 ] = 256'h00007fa0fffff631fffff631ffff8060ffff8060000009cf000009cf00007fa0;
    assign coff[305 ] = 256'h0000534fffff9ed2ffff9ed2ffffacb1ffffacb10000612e0000612e0000534f;
    assign coff[306 ] = 256'h00007228ffffc619ffffc619ffff8dd8ffff8dd8000039e7000039e700007228;
    assign coff[307 ] = 256'h000027c7ffff8656ffff8656ffffd839ffffd839000079aa000079aa000027c7;
    assign coff[308 ] = 256'h00007b42ffffdd7cffffdd7cffff84beffff84be000022840000228400007b42;
    assign coff[309 ] = 256'h00003ec0ffff9070ffff9070ffffc140ffffc14000006f9000006f9000003ec0;
    assign coff[310 ] = 256'h000064abffffb0f1ffffb0f1ffff9b55ffff9b5500004f0f00004f0f000064ab;
    assign coff[311 ] = 256'h00000f47ffff80eaffff80eafffff0b9fffff0b900007f1600007f1600000f47;
    assign coff[312 ] = 256'h00007e0cffffe9bbffffe9bbffff81f4ffff81f4000016450000164500007e0c;
    assign coff[313 ] = 256'h00004962ffff9720ffff9720ffffb69effffb69e000068e0000068e000004962;
    assign coff[314 ] = 256'h00006beeffffbb30ffffbb30ffff9412ffff9412000044d0000044d000006bee;
    assign coff[315 ] = 256'h00001ba9ffff8306ffff8306ffffe457ffffe45700007cfa00007cfa00001ba9;
    assign coff[316 ] = 256'h00007748ffffd191ffffd191ffff88b8ffff88b800002e6f00002e6f00007748;
    assign coff[317 ] = 256'h00003383ffff8ad3ffff8ad3ffffcc7dffffcc7d0000752d0000752d00003383;
    assign coff[318 ] = 256'h00005c6fffffa774ffffa774ffffa391ffffa3910000588c0000588c00005c6f;
    assign coff[319 ] = 256'h000002c0ffff8008ffff8008fffffd40fffffd4000007ff800007ff8000002c0;
    assign coff[320 ] = 256'h00007ffcfffffe09fffffe09ffff8004ffff8004000001f7000001f700007ffc;
    assign coff[321 ] = 256'h0000591cffffa41dffffa41dffffa6e4ffffa6e400005be300005be30000591c;
    assign coff[322 ] = 256'h0000757effffcd35ffffcd35ffff8a82ffff8a82000032cb000032cb0000757e;
    assign coff[323 ] = 256'h00002f2affff8902ffff8902ffffd0d6ffffd0d6000076fe000076fe00002f2a;
    assign coff[324 ] = 256'h00007d25ffffe51bffffe51bffff82dbffff82db00001ae500001ae500007d25;
    assign coff[325 ] = 256'h00004579ffff947effff947effffba87ffffba8700006b8200006b8200004579;
    assign coff[326 ] = 256'h00006953ffffb743ffffb743ffff96adffff96ad000048bd000048bd00006953;
    assign coff[327 ] = 256'h0000170bffff8217ffff8217ffffe8f5ffffe8f500007de900007de90000170b;
    assign coff[328 ] = 256'h00007f2dfffff180fffff180ffff80d3ffff80d300000e8000000e8000007f2d;
    assign coff[329 ] = 256'h00004fadffff9bd2ffff9bd2ffffb053ffffb0530000642e0000642e00004fad;
    assign coff[330 ] = 256'h00006ff2ffffc1f0ffffc1f0ffff900effff900e00003e1000003e1000006ff2;
    assign coff[331 ] = 256'h00002346ffff84f5ffff84f5ffffdcbaffffdcba00007b0b00007b0b00002346;
    assign coff[332 ] = 256'h000079e7ffffd8f8ffffd8f8ffff8619ffff86190000270800002708000079e7;
    assign coff[333 ] = 256'h00003a9affff8e34ffff8e34ffffc566ffffc566000071cc000071cc00003a9a;
    assign coff[334 ] = 256'h000061b0ffffad4affffad4affff9e50ffff9e50000052b6000052b6000061b0;
    assign coff[335 ] = 256'h00000a97ffff8070ffff8070fffff569fffff56900007f9000007f9000000a97;
    assign coff[336 ] = 256'h00007fbcfffff7c2fffff7c2ffff8044ffff80440000083e0000083e00007fbc;
    assign coff[337 ] = 256'h0000547fffff9fdaffff9fdaffffab81ffffab8100006026000060260000547f;
    assign coff[338 ] = 256'h000072dcffffc781ffffc781ffff8d24ffff8d240000387f0000387f000072dc;
    assign coff[339 ] = 256'h00002945ffff86d6ffff86d6ffffd6bbffffd6bb0000792a0000792a00002945;
    assign coff[340 ] = 256'h00007bacffffdeffffffdeffffff8454ffff8454000021010000210100007bac;
    assign coff[341 ] = 256'h0000401dffff9137ffff9137ffffbfe3ffffbfe300006ec900006ec90000401d;
    assign coff[342 ] = 256'h000065a1ffffb22fffffb22fffff9a5fffff9a5f00004dd100004dd1000065a1;
    assign coff[343 ] = 256'h000010d6ffff811dffff811dffffef2affffef2a00007ee300007ee3000010d6;
    assign coff[344 ] = 256'h00007e50ffffeb47ffffeb47ffff81b0ffff81b0000014b9000014b900007e50;
    assign coff[345 ] = 256'h00004aaaffff9808ffff9808ffffb556ffffb556000067f8000067f800004aaa;
    assign coff[346 ] = 256'h00006cc4ffffbc85ffffbc85ffff933cffff933c0000437b0000437b00006cc4;
    assign coff[347 ] = 256'h00001d31ffff8360ffff8360ffffe2cfffffe2cf00007ca000007ca000001d31;
    assign coff[348 ] = 256'h000077d8ffffd309ffffd309ffff8828ffff882800002cf700002cf7000077d8;
    assign coff[349 ] = 256'h000034f2ffff8b77ffff8b77ffffcb0effffcb0e0000748900007489000034f2;
    assign coff[350 ] = 256'h00005d83ffffa899ffffa899ffffa27dffffa27d000057670000576700005d83;
    assign coff[351 ] = 256'h00000452ffff8013ffff8013fffffbaefffffbae00007fed00007fed00000452;
    assign coff[352 ] = 256'h00007fe6fffffae5fffffae5ffff801affff801a0000051b0000051b00007fe6;
    assign coff[353 ] = 256'h000056d4ffffa1f4ffffa1f4ffffa92cffffa92c00005e0c00005e0c000056d4;
    assign coff[354 ] = 256'h00007436ffffca57ffffca57ffff8bcaffff8bca000035a9000035a900007436;
    assign coff[355 ] = 256'h00002c3bffff87e2ffff87e2ffffd3c5ffffd3c50000781e0000781e00002c3b;
    assign coff[356 ] = 256'h00007c72ffffe20bffffe20bffff838effff838e00001df500001df500007c72;
    assign coff[357 ] = 256'h000042d0ffff92d2ffff92d2ffffbd30ffffbd3000006d2e00006d2e000042d0;
    assign coff[358 ] = 256'h00006782ffffb4b3ffffb4b3ffff987effff987e00004b4d00004b4d00006782;
    assign coff[359 ] = 256'h000013f2ffff8190ffff8190ffffec0effffec0e00007e7000007e70000013f2;
    assign coff[360 ] = 256'h00007ec8ffffee62ffffee62ffff8138ffff81380000119e0000119e00007ec8;
    assign coff[361 ] = 256'h00004d31ffff99e5ffff99e5ffffb2cfffffb2cf0000661b0000661b00004d31;
    assign coff[362 ] = 256'h00006e64ffffbf35ffffbf35ffff919cffff919c000040cb000040cb00006e64;
    assign coff[363 ] = 256'h0000203effff8421ffff8421ffffdfc2ffffdfc200007bdf00007bdf0000203e;
    assign coff[364 ] = 256'h000078e9ffffd5fdffffd5fdffff8717ffff871700002a0300002a03000078e9;
    assign coff[365 ] = 256'h000037caffff8cccffff8cccffffc836ffffc8360000733400007334000037ca;
    assign coff[366 ] = 256'h00005fa1ffffaaebffffaaebffffa05fffffa05f000055150000551500005fa1;
    assign coff[367 ] = 256'h00000775ffff8038ffff8038fffff88bfffff88b00007fc800007fc800000775;
    assign coff[368 ] = 256'h00007f7efffff4a0fffff4a0ffff8082ffff808200000b6000000b6000007f7e;
    assign coff[369 ] = 256'h0000521cffff9dceffff9dceffffade4ffffade400006232000062320000521c;
    assign coff[370 ] = 256'h00007170ffffc4b4ffffc4b4ffff8e90ffff8e9000003b4c00003b4c00007170;
    assign coff[371 ] = 256'h00002648ffff85dcffff85dcffffd9b8ffffd9b800007a2400007a2400002648;
    assign coff[372 ] = 256'h00007ad3ffffdbf9ffffdbf9ffff852dffff852d000024070000240700007ad3;
    assign coff[373 ] = 256'h00003d60ffff8fadffff8fadffffc2a0ffffc2a0000070530000705300003d60;
    assign coff[374 ] = 256'h000063b0ffffafb6ffffafb6ffff9c50ffff9c500000504a0000504a000063b0;
    assign coff[375 ] = 256'h00000db8ffff80bdffff80bdfffff248fffff24800007f4300007f4300000db8;
    assign coff[376 ] = 256'h00007dc4ffffe82fffffe82fffff823cffff823c000017d1000017d100007dc4;
    assign coff[377 ] = 256'h00004817ffff963bffff963bffffb7e9ffffb7e9000069c5000069c500004817;
    assign coff[378 ] = 256'h00006b14ffffb9dfffffb9dfffff94ecffff94ec000046210000462100006b14;
    assign coff[379 ] = 256'h00001a20ffff82b2ffff82b2ffffe5e0ffffe5e000007d4e00007d4e00001a20;
    assign coff[380 ] = 256'h000076b4ffffd01bffffd01bffff894cffff894c00002fe500002fe5000076b4;
    assign coff[381 ] = 256'h00003212ffff8a33ffff8a33ffffcdeeffffcdee000075cd000075cd00003212;
    assign coff[382 ] = 256'h00005b57ffffa654ffffa654ffffa4a9ffffa4a9000059ac000059ac00005b57;
    assign coff[383 ] = 256'h0000012effff8001ffff8001fffffed2fffffed200007fff00007fff0000012e;
    assign coff[384 ] = 256'h00007ffffffffed2fffffed2ffff8001ffff80010000012e0000012e00007fff;
    assign coff[385 ] = 256'h000059acffffa4a9ffffa4a9ffffa654ffffa65400005b5700005b57000059ac;
    assign coff[386 ] = 256'h000075cdffffcdeeffffcdeeffff8a33ffff8a330000321200003212000075cd;
    assign coff[387 ] = 256'h00002fe5ffff894cffff894cffffd01bffffd01b000076b4000076b400002fe5;
    assign coff[388 ] = 256'h00007d4effffe5e0ffffe5e0ffff82b2ffff82b200001a2000001a2000007d4e;
    assign coff[389 ] = 256'h00004621ffff94ecffff94ecffffb9dfffffb9df00006b1400006b1400004621;
    assign coff[390 ] = 256'h000069c5ffffb7e9ffffb7e9ffff963bffff963b0000481700004817000069c5;
    assign coff[391 ] = 256'h000017d1ffff823cffff823cffffe82fffffe82f00007dc400007dc4000017d1;
    assign coff[392 ] = 256'h00007f43fffff248fffff248ffff80bdffff80bd00000db800000db800007f43;
    assign coff[393 ] = 256'h0000504affff9c50ffff9c50ffffafb6ffffafb6000063b0000063b00000504a;
    assign coff[394 ] = 256'h00007053ffffc2a0ffffc2a0ffff8fadffff8fad00003d6000003d6000007053;
    assign coff[395 ] = 256'h00002407ffff852dffff852dffffdbf9ffffdbf900007ad300007ad300002407;
    assign coff[396 ] = 256'h00007a24ffffd9b8ffffd9b8ffff85dcffff85dc000026480000264800007a24;
    assign coff[397 ] = 256'h00003b4cffff8e90ffff8e90ffffc4b4ffffc4b4000071700000717000003b4c;
    assign coff[398 ] = 256'h00006232ffffade4ffffade4ffff9dceffff9dce0000521c0000521c00006232;
    assign coff[399 ] = 256'h00000b60ffff8082ffff8082fffff4a0fffff4a000007f7e00007f7e00000b60;
    assign coff[400 ] = 256'h00007fc8fffff88bfffff88bffff8038ffff8038000007750000077500007fc8;
    assign coff[401 ] = 256'h00005515ffffa05fffffa05fffffaaebffffaaeb00005fa100005fa100005515;
    assign coff[402 ] = 256'h00007334ffffc836ffffc836ffff8cccffff8ccc000037ca000037ca00007334;
    assign coff[403 ] = 256'h00002a03ffff8717ffff8717ffffd5fdffffd5fd000078e9000078e900002a03;
    assign coff[404 ] = 256'h00007bdfffffdfc2ffffdfc2ffff8421ffff84210000203e0000203e00007bdf;
    assign coff[405 ] = 256'h000040cbffff919cffff919cffffbf35ffffbf3500006e6400006e64000040cb;
    assign coff[406 ] = 256'h0000661bffffb2cfffffb2cfffff99e5ffff99e500004d3100004d310000661b;
    assign coff[407 ] = 256'h0000119effff8138ffff8138ffffee62ffffee6200007ec800007ec80000119e;
    assign coff[408 ] = 256'h00007e70ffffec0effffec0effff8190ffff8190000013f2000013f200007e70;
    assign coff[409 ] = 256'h00004b4dffff987effff987effffb4b3ffffb4b3000067820000678200004b4d;
    assign coff[410 ] = 256'h00006d2effffbd30ffffbd30ffff92d2ffff92d2000042d0000042d000006d2e;
    assign coff[411 ] = 256'h00001df5ffff838effff838effffe20bffffe20b00007c7200007c7200001df5;
    assign coff[412 ] = 256'h0000781effffd3c5ffffd3c5ffff87e2ffff87e200002c3b00002c3b0000781e;
    assign coff[413 ] = 256'h000035a9ffff8bcaffff8bcaffffca57ffffca570000743600007436000035a9;
    assign coff[414 ] = 256'h00005e0cffffa92cffffa92cffffa1f4ffffa1f4000056d4000056d400005e0c;
    assign coff[415 ] = 256'h0000051bffff801affff801afffffae5fffffae500007fe600007fe60000051b;
    assign coff[416 ] = 256'h00007fedfffffbaefffffbaeffff8013ffff8013000004520000045200007fed;
    assign coff[417 ] = 256'h00005767ffffa27dffffa27dffffa899ffffa89900005d8300005d8300005767;
    assign coff[418 ] = 256'h00007489ffffcb0effffcb0effff8b77ffff8b77000034f2000034f200007489;
    assign coff[419 ] = 256'h00002cf7ffff8828ffff8828ffffd309ffffd309000077d8000077d800002cf7;
    assign coff[420 ] = 256'h00007ca0ffffe2cfffffe2cfffff8360ffff836000001d3100001d3100007ca0;
    assign coff[421 ] = 256'h0000437bffff933cffff933cffffbc85ffffbc8500006cc400006cc40000437b;
    assign coff[422 ] = 256'h000067f8ffffb556ffffb556ffff9808ffff980800004aaa00004aaa000067f8;
    assign coff[423 ] = 256'h000014b9ffff81b0ffff81b0ffffeb47ffffeb4700007e5000007e50000014b9;
    assign coff[424 ] = 256'h00007ee3ffffef2affffef2affff811dffff811d000010d6000010d600007ee3;
    assign coff[425 ] = 256'h00004dd1ffff9a5fffff9a5fffffb22fffffb22f000065a1000065a100004dd1;
    assign coff[426 ] = 256'h00006ec9ffffbfe3ffffbfe3ffff9137ffff91370000401d0000401d00006ec9;
    assign coff[427 ] = 256'h00002101ffff8454ffff8454ffffdeffffffdeff00007bac00007bac00002101;
    assign coff[428 ] = 256'h0000792affffd6bbffffd6bbffff86d6ffff86d600002945000029450000792a;
    assign coff[429 ] = 256'h0000387fffff8d24ffff8d24ffffc781ffffc781000072dc000072dc0000387f;
    assign coff[430 ] = 256'h00006026ffffab81ffffab81ffff9fdaffff9fda0000547f0000547f00006026;
    assign coff[431 ] = 256'h0000083effff8044ffff8044fffff7c2fffff7c200007fbc00007fbc0000083e;
    assign coff[432 ] = 256'h00007f90fffff569fffff569ffff8070ffff807000000a9700000a9700007f90;
    assign coff[433 ] = 256'h000052b6ffff9e50ffff9e50ffffad4affffad4a000061b0000061b0000052b6;
    assign coff[434 ] = 256'h000071ccffffc566ffffc566ffff8e34ffff8e3400003a9a00003a9a000071cc;
    assign coff[435 ] = 256'h00002708ffff8619ffff8619ffffd8f8ffffd8f8000079e7000079e700002708;
    assign coff[436 ] = 256'h00007b0bffffdcbaffffdcbaffff84f5ffff84f5000023460000234600007b0b;
    assign coff[437 ] = 256'h00003e10ffff900effff900effffc1f0ffffc1f000006ff200006ff200003e10;
    assign coff[438 ] = 256'h0000642effffb053ffffb053ffff9bd2ffff9bd200004fad00004fad0000642e;
    assign coff[439 ] = 256'h00000e80ffff80d3ffff80d3fffff180fffff18000007f2d00007f2d00000e80;
    assign coff[440 ] = 256'h00007de9ffffe8f5ffffe8f5ffff8217ffff82170000170b0000170b00007de9;
    assign coff[441 ] = 256'h000048bdffff96adffff96adffffb743ffffb7430000695300006953000048bd;
    assign coff[442 ] = 256'h00006b82ffffba87ffffba87ffff947effff947e000045790000457900006b82;
    assign coff[443 ] = 256'h00001ae5ffff82dbffff82dbffffe51bffffe51b00007d2500007d2500001ae5;
    assign coff[444 ] = 256'h000076feffffd0d6ffffd0d6ffff8902ffff890200002f2a00002f2a000076fe;
    assign coff[445 ] = 256'h000032cbffff8a82ffff8a82ffffcd35ffffcd350000757e0000757e000032cb;
    assign coff[446 ] = 256'h00005be3ffffa6e4ffffa6e4ffffa41dffffa41d0000591c0000591c00005be3;
    assign coff[447 ] = 256'h000001f7ffff8004ffff8004fffffe09fffffe0900007ffc00007ffc000001f7;
    assign coff[448 ] = 256'h00007ff8fffffd40fffffd40ffff8008ffff8008000002c0000002c000007ff8;
    assign coff[449 ] = 256'h0000588cffffa391ffffa391ffffa774ffffa77400005c6f00005c6f0000588c;
    assign coff[450 ] = 256'h0000752dffffcc7dffffcc7dffff8ad3ffff8ad300003383000033830000752d;
    assign coff[451 ] = 256'h00002e6fffff88b8ffff88b8ffffd191ffffd191000077480000774800002e6f;
    assign coff[452 ] = 256'h00007cfaffffe457ffffe457ffff8306ffff830600001ba900001ba900007cfa;
    assign coff[453 ] = 256'h000044d0ffff9412ffff9412ffffbb30ffffbb3000006bee00006bee000044d0;
    assign coff[454 ] = 256'h000068e0ffffb69effffb69effff9720ffff97200000496200004962000068e0;
    assign coff[455 ] = 256'h00001645ffff81f4ffff81f4ffffe9bbffffe9bb00007e0c00007e0c00001645;
    assign coff[456 ] = 256'h00007f16fffff0b9fffff0b9ffff80eaffff80ea00000f4700000f4700007f16;
    assign coff[457 ] = 256'h00004f0fffff9b55ffff9b55ffffb0f1ffffb0f1000064ab000064ab00004f0f;
    assign coff[458 ] = 256'h00006f90ffffc140ffffc140ffff9070ffff907000003ec000003ec000006f90;
    assign coff[459 ] = 256'h00002284ffff84beffff84beffffdd7cffffdd7c00007b4200007b4200002284;
    assign coff[460 ] = 256'h000079aaffffd839ffffd839ffff8656ffff8656000027c7000027c7000079aa;
    assign coff[461 ] = 256'h000039e7ffff8dd8ffff8dd8ffffc619ffffc6190000722800007228000039e7;
    assign coff[462 ] = 256'h0000612effffacb1ffffacb1ffff9ed2ffff9ed20000534f0000534f0000612e;
    assign coff[463 ] = 256'h000009cfffff8060ffff8060fffff631fffff63100007fa000007fa0000009cf;
    assign coff[464 ] = 256'h00007faefffff6fafffff6faffff8052ffff8052000009060000090600007fae;
    assign coff[465 ] = 256'h000053e7ffff9f56ffff9f56ffffac19ffffac19000060aa000060aa000053e7;
    assign coff[466 ] = 256'h00007282ffffc6cdffffc6cdffff8d7effff8d7e000039330000393300007282;
    assign coff[467 ] = 256'h00002886ffff8696ffff8696ffffd77affffd77a0000796a0000796a00002886;
    assign coff[468 ] = 256'h00007b78ffffde3dffffde3dffff8488ffff8488000021c3000021c300007b78;
    assign coff[469 ] = 256'h00003f6fffff90d3ffff90d3ffffc091ffffc09100006f2d00006f2d00003f6f;
    assign coff[470 ] = 256'h00006526ffffb18fffffb18fffff9adaffff9ada00004e7100004e7100006526;
    assign coff[471 ] = 256'h0000100fffff8103ffff8103ffffeff1ffffeff100007efd00007efd0000100f;
    assign coff[472 ] = 256'h00007e2fffffea81ffffea81ffff81d1ffff81d10000157f0000157f00007e2f;
    assign coff[473 ] = 256'h00004a06ffff9793ffff9793ffffb5faffffb5fa0000686d0000686d00004a06;
    assign coff[474 ] = 256'h00006c5affffbbdaffffbbdaffff93a6ffff93a6000044260000442600006c5a;
    assign coff[475 ] = 256'h00001c6effff8332ffff8332ffffe392ffffe39200007cce00007cce00001c6e;
    assign coff[476 ] = 256'h00007790ffffd24dffffd24dffff8870ffff887000002db300002db300007790;
    assign coff[477 ] = 256'h0000343bffff8b24ffff8b24ffffcbc5ffffcbc5000074dc000074dc0000343b;
    assign coff[478 ] = 256'h00005cf9ffffa806ffffa806ffffa307ffffa307000057fa000057fa00005cf9;
    assign coff[479 ] = 256'h00000389ffff800cffff800cfffffc77fffffc7700007ff400007ff400000389;
    assign coff[480 ] = 256'h00007fddfffffa1dfffffa1dffff8023ffff8023000005e3000005e300007fdd;
    assign coff[481 ] = 256'h00005640ffffa16cffffa16cffffa9c0ffffa9c000005e9400005e9400005640;
    assign coff[482 ] = 256'h000073e1ffffc9a1ffffc9a1ffff8c1fffff8c1f0000365f0000365f000073e1;
    assign coff[483 ] = 256'h00002b7effff879dffff879dffffd482ffffd482000078630000786300002b7e;
    assign coff[484 ] = 256'h00007c42ffffe148ffffe148ffff83beffff83be00001eb800001eb800007c42;
    assign coff[485 ] = 256'h00004224ffff926affff926affffbddcffffbddc00006d9600006d9600004224;
    assign coff[486 ] = 256'h0000670bffffb411ffffb411ffff98f5ffff98f500004bef00004bef0000670b;
    assign coff[487 ] = 256'h0000132bffff8172ffff8172ffffecd5ffffecd500007e8e00007e8e0000132b;
    assign coff[488 ] = 256'h00007eacffffed9bffffed9bffff8154ffff8154000012650000126500007eac;
    assign coff[489 ] = 256'h00004c91ffff996dffff996dffffb36fffffb36f000066930000669300004c91;
    assign coff[490 ] = 256'h00006dfeffffbe88ffffbe88ffff9202ffff9202000041780000417800006dfe;
    assign coff[491 ] = 256'h00001f7bffff83efffff83efffffe085ffffe08500007c1100007c1100001f7b;
    assign coff[492 ] = 256'h000078a6ffffd53fffffd53fffff875affff875a00002ac100002ac1000078a6;
    assign coff[493 ] = 256'h00003715ffff8c75ffff8c75ffffc8ebffffc8eb0000738b0000738b00003715;
    assign coff[494 ] = 256'h00005f1bffffaa55ffffaa55ffffa0e5ffffa0e5000055ab000055ab00005f1b;
    assign coff[495 ] = 256'h000006acffff802dffff802dfffff954fffff95400007fd300007fd3000006ac;
    assign coff[496 ] = 256'h00007f6cfffff3d8fffff3d8ffff8094ffff809400000c2800000c2800007f6c;
    assign coff[497 ] = 256'h00005181ffff9d4effff9d4effffae7fffffae7f000062b2000062b200005181;
    assign coff[498 ] = 256'h00007112ffffc402ffffc402ffff8eeeffff8eee00003bfe00003bfe00007112;
    assign coff[499 ] = 256'h00002588ffff85a0ffff85a0ffffda78ffffda7800007a6000007a6000002588;
    assign coff[500 ] = 256'h00007a9affffdb38ffffdb38ffff8566ffff8566000024c8000024c800007a9a;
    assign coff[501 ] = 256'h00003cafffff8f4dffff8f4dffffc351ffffc351000070b3000070b300003caf;
    assign coff[502 ] = 256'h00006332ffffaf1affffaf1affff9cceffff9cce000050e6000050e600006332;
    assign coff[503 ] = 256'h00000cf0ffff80a8ffff80a8fffff310fffff31000007f5800007f5800000cf0;
    assign coff[504 ] = 256'h00007d9effffe76affffe76affff8262ffff8262000018960000189600007d9e;
    assign coff[505 ] = 256'h00004770ffff95caffff95caffffb890ffffb89000006a3600006a3600004770;
    assign coff[506 ] = 256'h00006aa5ffffb937ffffb937ffff955bffff955b000046c9000046c900006aa5;
    assign coff[507 ] = 256'h0000195bffff8289ffff8289ffffe6a5ffffe6a500007d7700007d770000195b;
    assign coff[508 ] = 256'h00007668ffffcf61ffffcf61ffff8998ffff89980000309f0000309f00007668;
    assign coff[509 ] = 256'h00003159ffff89e5ffff89e5ffffcea7ffffcea70000761b0000761b00003159;
    assign coff[510 ] = 256'h00005ac9ffffa5c5ffffa5c5ffffa537ffffa53700005a3b00005a3b00005ac9;
    assign coff[511 ] = 256'h00000065ffff8001ffff8001ffffff9bffffff9b00007fff00007fff00000065;
    assign coff[512 ] = 256'h00007fffffffffceffffffceffff8001ffff8001000000320000003200007fff;
    assign coff[513 ] = 256'h00005a5fffffa55affffa55affffa5a1ffffa5a100005aa600005aa600005a5f;
    assign coff[514 ] = 256'h0000762effffced6ffffced6ffff89d2ffff89d20000312a0000312a0000762e;
    assign coff[515 ] = 256'h000030cdffff89abffff89abffffcf33ffffcf330000765500007655000030cd;
    assign coff[516 ] = 256'h00007d81ffffe6d6ffffe6d6ffff827fffff827f0000192a0000192a00007d81;
    assign coff[517 ] = 256'h000046f3ffff9577ffff9577ffffb90dffffb90d00006a8900006a89000046f3;
    assign coff[518 ] = 256'h00006a52ffffb8b9ffffb8b9ffff95aeffff95ae000047470000474700006a52;
    assign coff[519 ] = 256'h000018c7ffff826cffff826cffffe739ffffe73900007d9400007d94000018c7;
    assign coff[520 ] = 256'h00007f5dfffff342fffff342ffff80a3ffff80a300000cbe00000cbe00007f5d;
    assign coff[521 ] = 256'h0000510dffff9ceeffff9ceeffffaef3ffffaef300006312000063120000510d;
    assign coff[522 ] = 256'h000070cbffffc37dffffc37dffff8f35ffff8f3500003c8300003c83000070cb;
    assign coff[523 ] = 256'h000024f8ffff8574ffff8574ffffdb08ffffdb0800007a8c00007a8c000024f8;
    assign coff[524 ] = 256'h00007a6effffdaa8ffffdaa8ffff8592ffff8592000025580000255800007a6e;
    assign coff[525 ] = 256'h00003c2affff8f06ffff8f06ffffc3d6ffffc3d6000070fa000070fa00003c2a;
    assign coff[526 ] = 256'h000062d2ffffaea5ffffaea5ffff9d2effff9d2e0000515b0000515b000062d2;
    assign coff[527 ] = 256'h00000c5affff8099ffff8099fffff3a6fffff3a600007f6700007f6700000c5a;
    assign coff[528 ] = 256'h00007fd6fffff986fffff986ffff802affff802a0000067a0000067a00007fd6;
    assign coff[529 ] = 256'h000055d0ffffa107ffffa107ffffaa30ffffaa3000005ef900005ef9000055d0;
    assign coff[530 ] = 256'h000073a0ffffc918ffffc918ffff8c60ffff8c60000036e8000036e8000073a0;
    assign coff[531 ] = 256'h00002af0ffff876bffff876bffffd510ffffd510000078950000789500002af0;
    assign coff[532 ] = 256'h00007c1effffe0b5ffffe0b5ffff83e2ffff83e200001f4b00001f4b00007c1e;
    assign coff[533 ] = 256'h000041a3ffff921cffff921cffffbe5dffffbe5d00006de400006de4000041a3;
    assign coff[534 ] = 256'h000066b2ffffb398ffffb398ffff994effff994e00004c6800004c68000066b2;
    assign coff[535 ] = 256'h00001296ffff815bffff815bffffed6affffed6a00007ea500007ea500001296;
    assign coff[536 ] = 256'h00007e96ffffed06ffffed06ffff816affff816a000012fa000012fa00007e96;
    assign coff[537 ] = 256'h00004c17ffff9913ffff9913ffffb3e9ffffb3e9000066ed000066ed00004c17;
    assign coff[538 ] = 256'h00006db0ffffbe07ffffbe07ffff9250ffff9250000041f9000041f900006db0;
    assign coff[539 ] = 256'h00001ee9ffff83caffff83caffffe117ffffe11700007c3600007c3600001ee9;
    assign coff[540 ] = 256'h00007874ffffd4b1ffffd4b1ffff878cffff878c00002b4f00002b4f00007874;
    assign coff[541 ] = 256'h0000368dffff8c35ffff8c35ffffc973ffffc973000073cb000073cb0000368d;
    assign coff[542 ] = 256'h00005eb6ffffa9e5ffffa9e5ffffa14affffa14a0000561b0000561b00005eb6;
    assign coff[543 ] = 256'h00000616ffff8025ffff8025fffff9eafffff9ea00007fdb00007fdb00000616;
    assign coff[544 ] = 256'h00007ff5fffffcaafffffcaaffff800bffff800b000003560000035600007ff5;
    assign coff[545 ] = 256'h0000581effffa329ffffa329ffffa7e2ffffa7e200005cd700005cd70000581e;
    assign coff[546 ] = 256'h000074f0ffffcbf3ffffcbf3ffff8b10ffff8b100000340d0000340d000074f0;
    assign coff[547 ] = 256'h00002de2ffff8882ffff8882ffffd21effffd21e0000777e0000777e00002de2;
    assign coff[548 ] = 256'h00007cd9ffffe3c3ffffe3c3ffff8327ffff832700001c3d00001c3d00007cd9;
    assign coff[549 ] = 256'h00004450ffff93c1ffff93c1ffffbbb0ffffbbb000006c3f00006c3f00004450;
    assign coff[550 ] = 256'h0000688affffb623ffffb623ffff9776ffff9776000049dd000049dd0000688a;
    assign coff[551 ] = 256'h000015b1ffff81daffff81daffffea4fffffea4f00007e2600007e26000015b1;
    assign coff[552 ] = 256'h00007f03fffff023fffff023ffff80fdffff80fd00000fdd00000fdd00007f03;
    assign coff[553 ] = 256'h00004e98ffff9af9ffff9af9ffffb168ffffb168000065070000650700004e98;
    assign coff[554 ] = 256'h00006f46ffffc0bdffffc0bdffff90baffff90ba00003f4300003f4300006f46;
    assign coff[555 ] = 256'h000021f3ffff8496ffff8496ffffde0dffffde0d00007b6a00007b6a000021f3;
    assign coff[556 ] = 256'h0000797affffd7aaffffd7aaffff8686ffff868600002856000028560000797a;
    assign coff[557 ] = 256'h00003960ffff8d94ffff8d94ffffc6a0ffffc6a00000726c0000726c00003960;
    assign coff[558 ] = 256'h000060cbffffac3fffffac3fffff9f35ffff9f35000053c1000053c1000060cb;
    assign coff[559 ] = 256'h00000938ffff8055ffff8055fffff6c8fffff6c800007fab00007fab00000938;
    assign coff[560 ] = 256'h00007fa3fffff663fffff663ffff805dffff805d0000099d0000099d00007fa3;
    assign coff[561 ] = 256'h00005375ffff9ef3ffff9ef3ffffac8bffffac8b0000610d0000610d00005375;
    assign coff[562 ] = 256'h0000723fffffc646ffffc646ffff8dc1ffff8dc1000039ba000039ba0000723f;
    assign coff[563 ] = 256'h000027f7ffff8666ffff8666ffffd809ffffd8090000799a0000799a000027f7;
    assign coff[564 ] = 256'h00007b50ffffddacffffddacffff84b0ffff84b0000022540000225400007b50;
    assign coff[565 ] = 256'h00003eecffff9088ffff9088ffffc114ffffc11400006f7800006f7800003eec;
    assign coff[566 ] = 256'h000064caffffb118ffffb118ffff9b36ffff9b3600004ee800004ee8000064ca;
    assign coff[567 ] = 256'h00000f79ffff80f0ffff80f0fffff087fffff08700007f1000007f1000000f79;
    assign coff[568 ] = 256'h00007e15ffffe9ecffffe9ecffff81ebffff81eb000016140000161400007e15;
    assign coff[569 ] = 256'h0000498bffff973cffff973cffffb675ffffb675000068c4000068c40000498b;
    assign coff[570 ] = 256'h00006c09ffffbb5bffffbb5bffff93f7ffff93f7000044a5000044a500006c09;
    assign coff[571 ] = 256'h00001bdaffff8311ffff8311ffffe426ffffe42600007cef00007cef00001bda;
    assign coff[572 ] = 256'h0000775affffd1c0ffffd1c0ffff88a6ffff88a600002e4000002e400000775a;
    assign coff[573 ] = 256'h000033b1ffff8ae7ffff8ae7ffffcc4fffffcc4f0000751900007519000033b1;
    assign coff[574 ] = 256'h00005c91ffffa799ffffa799ffffa36fffffa36f000058670000586700005c91;
    assign coff[575 ] = 256'h000002f2ffff8009ffff8009fffffd0efffffd0e00007ff700007ff7000002f2;
    assign coff[576 ] = 256'h00007ffdfffffe3cfffffe3cffff8003ffff8003000001c4000001c400007ffd;
    assign coff[577 ] = 256'h00005940ffffa440ffffa440ffffa6c0ffffa6c000005bc000005bc000005940;
    assign coff[578 ] = 256'h00007592ffffcd63ffffcd63ffff8a6effff8a6e0000329d0000329d00007592;
    assign coff[579 ] = 256'h00002f59ffff8914ffff8914ffffd0a7ffffd0a7000076ec000076ec00002f59;
    assign coff[580 ] = 256'h00007d2fffffe54cffffe54cffff82d1ffff82d100001ab400001ab400007d2f;
    assign coff[581 ] = 256'h000045a3ffff949affff949affffba5dffffba5d00006b6600006b66000045a3;
    assign coff[582 ] = 256'h00006970ffffb76dffffb76dffff9690ffff9690000048930000489300006970;
    assign coff[583 ] = 256'h0000173cffff8220ffff8220ffffe8c4ffffe8c400007de000007de00000173c;
    assign coff[584 ] = 256'h00007f33fffff1b2fffff1b2ffff80cdffff80cd00000e4e00000e4e00007f33;
    assign coff[585 ] = 256'h00004fd4ffff9bf1ffff9bf1ffffb02cffffb02c0000640f0000640f00004fd4;
    assign coff[586 ] = 256'h0000700bffffc21cffffc21cffff8ff5ffff8ff500003de400003de40000700b;
    assign coff[587 ] = 256'h00002376ffff8503ffff8503ffffdc8affffdc8a00007afd00007afd00002376;
    assign coff[588 ] = 256'h000079f7ffffd928ffffd928ffff8609ffff8609000026d8000026d8000079f7;
    assign coff[589 ] = 256'h00003ac6ffff8e4bffff8e4bffffc53affffc53a000071b5000071b500003ac6;
    assign coff[590 ] = 256'h000061d1ffffad70ffffad70ffff9e2fffff9e2f0000529000005290000061d1;
    assign coff[591 ] = 256'h00000ac9ffff8075ffff8075fffff537fffff53700007f8b00007f8b00000ac9;
    assign coff[592 ] = 256'h00007fbffffff7f4fffff7f4ffff8041ffff80410000080c0000080c00007fbf;
    assign coff[593 ] = 256'h000054a4ffff9ffbffff9ffbffffab5cffffab5c0000600500006005000054a4;
    assign coff[594 ] = 256'h000072f2ffffc7aeffffc7aeffff8d0effff8d0e0000385200003852000072f2;
    assign coff[595 ] = 256'h00002974ffff86e6ffff86e6ffffd68cffffd68c0000791a0000791a00002974;
    assign coff[596 ] = 256'h00007bb9ffffdf30ffffdf30ffff8447ffff8447000020d0000020d000007bb9;
    assign coff[597 ] = 256'h00004048ffff9150ffff9150ffffbfb8ffffbfb800006eb000006eb000004048;
    assign coff[598 ] = 256'h000065c0ffffb257ffffb257ffff9a40ffff9a4000004da900004da9000065c0;
    assign coff[599 ] = 256'h00001108ffff8123ffff8123ffffeef8ffffeef800007edd00007edd00001108;
    assign coff[600 ] = 256'h00007e58ffffeb79ffffeb79ffff81a8ffff81a8000014870000148700007e58;
    assign coff[601 ] = 256'h00004ad3ffff9826ffff9826ffffb52dffffb52d000067da000067da00004ad3;
    assign coff[602 ] = 256'h00006cdfffffbcafffffbcafffff9321ffff9321000043510000435100006cdf;
    assign coff[603 ] = 256'h00001d62ffff836bffff836bffffe29effffe29e00007c9500007c9500001d62;
    assign coff[604 ] = 256'h000077e9ffffd338ffffd338ffff8817ffff881700002cc800002cc8000077e9;
    assign coff[605 ] = 256'h00003520ffff8b8bffff8b8bffffcae0ffffcae0000074750000747500003520;
    assign coff[606 ] = 256'h00005da5ffffa8bdffffa8bdffffa25bffffa25b000057430000574300005da5;
    assign coff[607 ] = 256'h00000484ffff8014ffff8014fffffb7cfffffb7c00007fec00007fec00000484;
    assign coff[608 ] = 256'h00007fe8fffffb18fffffb18ffff8018ffff8018000004e8000004e800007fe8;
    assign coff[609 ] = 256'h000056f9ffffa216ffffa216ffffa907ffffa90700005dea00005dea000056f9;
    assign coff[610 ] = 256'h0000744bffffca85ffffca85ffff8bb5ffff8bb50000357b0000357b0000744b;
    assign coff[611 ] = 256'h00002c6affff87f4ffff87f4ffffd396ffffd3960000780c0000780c00002c6a;
    assign coff[612 ] = 256'h00007c7effffe23cffffe23cffff8382ffff838200001dc400001dc400007c7e;
    assign coff[613 ] = 256'h000042fbffff92ecffff92ecffffbd05ffffbd0500006d1400006d14000042fb;
    assign coff[614 ] = 256'h000067a0ffffb4dcffffb4dcffff9860ffff986000004b2400004b24000067a0;
    assign coff[615 ] = 256'h00001424ffff8198ffff8198ffffebdcffffebdc00007e6800007e6800001424;
    assign coff[616 ] = 256'h00007ecfffffee94ffffee94ffff8131ffff81310000116c0000116c00007ecf;
    assign coff[617 ] = 256'h00004d59ffff9a04ffff9a04ffffb2a7ffffb2a7000065fc000065fc00004d59;
    assign coff[618 ] = 256'h00006e7dffffbf61ffffbf61ffff9183ffff91830000409f0000409f00006e7d;
    assign coff[619 ] = 256'h0000206fffff842dffff842dffffdf91ffffdf9100007bd300007bd30000206f;
    assign coff[620 ] = 256'h000078f9ffffd62dffffd62dffff8707ffff8707000029d3000029d3000078f9;
    assign coff[621 ] = 256'h000037f7ffff8ce2ffff8ce2ffffc809ffffc8090000731e0000731e000037f7;
    assign coff[622 ] = 256'h00005fc2ffffab10ffffab10ffffa03effffa03e000054f0000054f000005fc2;
    assign coff[623 ] = 256'h000007a7ffff803bffff803bfffff859fffff85900007fc500007fc5000007a7;
    assign coff[624 ] = 256'h00007f83fffff4d3fffff4d3ffff807dffff807d00000b2d00000b2d00007f83;
    assign coff[625 ] = 256'h00005243ffff9defffff9defffffadbdffffadbd000062110000621100005243;
    assign coff[626 ] = 256'h00007187ffffc4e0ffffc4e0ffff8e79ffff8e7900003b2000003b2000007187;
    assign coff[627 ] = 256'h00002678ffff85ebffff85ebffffd988ffffd98800007a1500007a1500002678;
    assign coff[628 ] = 256'h00007ae1ffffdc29ffffdc29ffff851fffff851f000023d7000023d700007ae1;
    assign coff[629 ] = 256'h00003d8cffff8fc5ffff8fc5ffffc274ffffc2740000703b0000703b00003d8c;
    assign coff[630 ] = 256'h000063d0ffffafddffffafddffff9c30ffff9c300000502300005023000063d0;
    assign coff[631 ] = 256'h00000deaffff80c2ffff80c2fffff216fffff21600007f3e00007f3e00000dea;
    assign coff[632 ] = 256'h00007dcdffffe861ffffe861ffff8233ffff82330000179f0000179f00007dcd;
    assign coff[633 ] = 256'h00004840ffff9657ffff9657ffffb7c0ffffb7c0000069a9000069a900004840;
    assign coff[634 ] = 256'h00006b30ffffba09ffffba09ffff94d0ffff94d0000045f7000045f700006b30;
    assign coff[635 ] = 256'h00001a51ffff82bcffff82bcffffe5afffffe5af00007d4400007d4400001a51;
    assign coff[636 ] = 256'h000076c7ffffd04affffd04affff8939ffff893900002fb600002fb6000076c7;
    assign coff[637 ] = 256'h00003240ffff8a47ffff8a47ffffcdc0ffffcdc0000075b9000075b900003240;
    assign coff[638 ] = 256'h00005b7affffa678ffffa678ffffa486ffffa486000059880000598800005b7a;
    assign coff[639 ] = 256'h00000160ffff8002ffff8002fffffea0fffffea000007ffe00007ffe00000160;
    assign coff[640 ] = 256'h00007fffffffff05ffffff05ffff8001ffff8001000000fb000000fb00007fff;
    assign coff[641 ] = 256'h000059d0ffffa4ccffffa4ccffffa630ffffa63000005b3400005b34000059d0;
    assign coff[642 ] = 256'h000075e1ffffce1cffffce1cffff8a1fffff8a1f000031e4000031e4000075e1;
    assign coff[643 ] = 256'h00003013ffff895fffff895fffffcfedffffcfed000076a1000076a100003013;
    assign coff[644 ] = 256'h00007d58ffffe611ffffe611ffff82a8ffff82a8000019ef000019ef00007d58;
    assign coff[645 ] = 256'h0000464bffff9508ffff9508ffffb9b5ffffb9b500006af800006af80000464b;
    assign coff[646 ] = 256'h000069e1ffffb813ffffb813ffff961fffff961f000047ed000047ed000069e1;
    assign coff[647 ] = 256'h00001802ffff8246ffff8246ffffe7feffffe7fe00007dba00007dba00001802;
    assign coff[648 ] = 256'h00007f49fffff27afffff27affff80b7ffff80b700000d8600000d8600007f49;
    assign coff[649 ] = 256'h00005071ffff9c6fffff9c6fffffaf8fffffaf8f000063910000639100005071;
    assign coff[650 ] = 256'h0000706bffffc2ccffffc2ccffff8f95ffff8f9500003d3400003d340000706b;
    assign coff[651 ] = 256'h00002437ffff853bffff853bffffdbc9ffffdbc900007ac500007ac500002437;
    assign coff[652 ] = 256'h00007a33ffffd9e8ffffd9e8ffff85cdffff85cd000026180000261800007a33;
    assign coff[653 ] = 256'h00003b79ffff8ea8ffff8ea8ffffc487ffffc487000071580000715800003b79;
    assign coff[654 ] = 256'h00006252ffffae0bffffae0bffff9daeffff9dae000051f5000051f500006252;
    assign coff[655 ] = 256'h00000b92ffff8086ffff8086fffff46efffff46e00007f7a00007f7a00000b92;
    assign coff[656 ] = 256'h00007fcbfffff8bdfffff8bdffff8035ffff8035000007430000074300007fcb;
    assign coff[657 ] = 256'h0000553bffffa080ffffa080ffffaac5ffffaac500005f8000005f800000553b;
    assign coff[658 ] = 256'h0000734affffc863ffffc863ffff8cb6ffff8cb60000379d0000379d0000734a;
    assign coff[659 ] = 256'h00002a32ffff8728ffff8728ffffd5ceffffd5ce000078d8000078d800002a32;
    assign coff[660 ] = 256'h00007becffffdff2ffffdff2ffff8414ffff84140000200e0000200e00007bec;
    assign coff[661 ] = 256'h000040f6ffff91b6ffff91b6ffffbf0affffbf0a00006e4a00006e4a000040f6;
    assign coff[662 ] = 256'h00006639ffffb2f7ffffb2f7ffff99c7ffff99c700004d0900004d0900006639;
    assign coff[663 ] = 256'h000011cfffff813fffff813fffffee31ffffee3100007ec100007ec1000011cf;
    assign coff[664 ] = 256'h00007e78ffffec3fffffec3fffff8188ffff8188000013c1000013c100007e78;
    assign coff[665 ] = 256'h00004b75ffff989cffff989cffffb48bffffb48b000067640000676400004b75;
    assign coff[666 ] = 256'h00006d48ffffbd5bffffbd5bffff92b8ffff92b8000042a5000042a500006d48;
    assign coff[667 ] = 256'h00001e26ffff839affff839affffe1daffffe1da00007c6600007c6600001e26;
    assign coff[668 ] = 256'h0000782fffffd3f4ffffd3f4ffff87d1ffff87d100002c0c00002c0c0000782f;
    assign coff[669 ] = 256'h000035d7ffff8bdfffff8bdfffffca29ffffca290000742100007421000035d7;
    assign coff[670 ] = 256'h00005e2effffa951ffffa951ffffa1d2ffffa1d2000056af000056af00005e2e;
    assign coff[671 ] = 256'h0000054dffff801cffff801cfffffab3fffffab300007fe400007fe40000054d;
    assign coff[672 ] = 256'h00007feffffffbe1fffffbe1ffff8011ffff80110000041f0000041f00007fef;
    assign coff[673 ] = 256'h0000578cffffa29fffffa29fffffa874ffffa87400005d6100005d610000578c;
    assign coff[674 ] = 256'h0000749effffcb3cffffcb3cffff8b62ffff8b62000034c4000034c40000749e;
    assign coff[675 ] = 256'h00002d26ffff883affff883affffd2daffffd2da000077c6000077c600002d26;
    assign coff[676 ] = 256'h00007cacffffe2ffffffe2ffffff8354ffff835400001d0100001d0100007cac;
    assign coff[677 ] = 256'h000043a6ffff9356ffff9356ffffbc5affffbc5a00006caa00006caa000043a6;
    assign coff[678 ] = 256'h00006815ffffb57fffffb57fffff97ebffff97eb00004a8100004a8100006815;
    assign coff[679 ] = 256'h000014eaffff81b8ffff81b8ffffeb16ffffeb1600007e4800007e48000014ea;
    assign coff[680 ] = 256'h00007eeaffffef5cffffef5cffff8116ffff8116000010a4000010a400007eea;
    assign coff[681 ] = 256'h00004df9ffff9a7effff9a7effffb207ffffb207000065820000658200004df9;
    assign coff[682 ] = 256'h00006ee2ffffc00fffffc00fffff911effff911e00003ff100003ff100006ee2;
    assign coff[683 ] = 256'h00002131ffff8461ffff8461ffffdecfffffdecf00007b9f00007b9f00002131;
    assign coff[684 ] = 256'h0000793affffd6ebffffd6ebffff86c6ffff86c600002915000029150000793a;
    assign coff[685 ] = 256'h000038acffff8d3bffff8d3bffffc754ffffc754000072c5000072c5000038ac;
    assign coff[686 ] = 256'h00006047ffffaba7ffffaba7ffff9fb9ffff9fb9000054590000545900006047;
    assign coff[687 ] = 256'h00000870ffff8047ffff8047fffff790fffff79000007fb900007fb900000870;
    assign coff[688 ] = 256'h00007f94fffff59bfffff59bffff806cffff806c00000a6500000a6500007f94;
    assign coff[689 ] = 256'h000052dcffff9e70ffff9e70ffffad24ffffad240000619000006190000052dc;
    assign coff[690 ] = 256'h000071e3ffffc593ffffc593ffff8e1dffff8e1d00003a6d00003a6d000071e3;
    assign coff[691 ] = 256'h00002738ffff8628ffff8628ffffd8c8ffffd8c8000079d8000079d800002738;
    assign coff[692 ] = 256'h00007b19ffffdceaffffdceaffff84e7ffff84e7000023160000231600007b19;
    assign coff[693 ] = 256'h00003e3cffff9026ffff9026ffffc1c4ffffc1c400006fda00006fda00003e3c;
    assign coff[694 ] = 256'h0000644dffffb07bffffb07bffff9bb3ffff9bb300004f8500004f850000644d;
    assign coff[695 ] = 256'h00000eb2ffff80d9ffff80d9fffff14efffff14e00007f2700007f2700000eb2;
    assign coff[696 ] = 256'h00007df2ffffe926ffffe926ffff820effff820e000016da000016da00007df2;
    assign coff[697 ] = 256'h000048e6ffff96c9ffff96c9ffffb71affffb71a0000693700006937000048e6;
    assign coff[698 ] = 256'h00006b9dffffbab1ffffbab1ffff9463ffff94630000454f0000454f00006b9d;
    assign coff[699 ] = 256'h00001b16ffff82e6ffff82e6ffffe4eaffffe4ea00007d1a00007d1a00001b16;
    assign coff[700 ] = 256'h00007711ffffd105ffffd105ffff88efffff88ef00002efb00002efb00007711;
    assign coff[701 ] = 256'h000032f9ffff8a96ffff8a96ffffcd07ffffcd070000756a0000756a000032f9;
    assign coff[702 ] = 256'h00005c06ffffa708ffffa708ffffa3faffffa3fa000058f8000058f800005c06;
    assign coff[703 ] = 256'h00000229ffff8005ffff8005fffffdd7fffffdd700007ffb00007ffb00000229;
    assign coff[704 ] = 256'h00007ff9fffffd73fffffd73ffff8007ffff80070000028d0000028d00007ff9;
    assign coff[705 ] = 256'h000058b0ffffa3b4ffffa3b4ffffa750ffffa75000005c4c00005c4c000058b0;
    assign coff[706 ] = 256'h00007542ffffccabffffccabffff8abeffff8abe000033550000335500007542;
    assign coff[707 ] = 256'h00002e9effff88caffff88caffffd162ffffd162000077360000773600002e9e;
    assign coff[708 ] = 256'h00007d05ffffe488ffffe488ffff82fbffff82fb00001b7800001b7800007d05;
    assign coff[709 ] = 256'h000044faffff942dffff942dffffbb06ffffbb0600006bd300006bd3000044fa;
    assign coff[710 ] = 256'h000068fdffffb6c7ffffb6c7ffff9703ffff97030000493900004939000068fd;
    assign coff[711 ] = 256'h00001677ffff81fdffff81fdffffe989ffffe98900007e0300007e0300001677;
    assign coff[712 ] = 256'h00007f1cfffff0ebfffff0ebffff80e4ffff80e400000f1500000f1500007f1c;
    assign coff[713 ] = 256'h00004f37ffff9b75ffff9b75ffffb0c9ffffb0c90000648b0000648b00004f37;
    assign coff[714 ] = 256'h00006fa9ffffc16cffffc16cffff9057ffff905700003e9400003e9400006fa9;
    assign coff[715 ] = 256'h000022b5ffff84ccffff84ccffffdd4bffffdd4b00007b3400007b34000022b5;
    assign coff[716 ] = 256'h000079b9ffffd869ffffd869ffff8647ffff86470000279700002797000079b9;
    assign coff[717 ] = 256'h00003a13ffff8defffff8defffffc5edffffc5ed000072110000721100003a13;
    assign coff[718 ] = 256'h0000614effffacd7ffffacd7ffff9eb2ffff9eb200005329000053290000614e;
    assign coff[719 ] = 256'h00000a01ffff8064ffff8064fffff5fffffff5ff00007f9c00007f9c00000a01;
    assign coff[720 ] = 256'h00007fb2fffff72cfffff72cffff804effff804e000008d4000008d400007fb2;
    assign coff[721 ] = 256'h0000540dffff9f77ffff9f77ffffabf3ffffabf300006089000060890000540d;
    assign coff[722 ] = 256'h00007299ffffc6faffffc6faffff8d67ffff8d67000039060000390600007299;
    assign coff[723 ] = 256'h000028b6ffff86a5ffff86a5ffffd74affffd74a0000795b0000795b000028b6;
    assign coff[724 ] = 256'h00007b85ffffde6effffde6effff847bffff847b000021920000219200007b85;
    assign coff[725 ] = 256'h00003f9affff90ecffff90ecffffc066ffffc06600006f1400006f1400003f9a;
    assign coff[726 ] = 256'h00006545ffffb1b7ffffb1b7ffff9abbffff9abb00004e4900004e4900006545;
    assign coff[727 ] = 256'h00001041ffff8109ffff8109ffffefbfffffefbf00007ef700007ef700001041;
    assign coff[728 ] = 256'h00007e37ffffeab3ffffeab3ffff81c9ffff81c90000154d0000154d00007e37;
    assign coff[729 ] = 256'h00004a2fffff97b0ffff97b0ffffb5d1ffffb5d1000068500000685000004a2f;
    assign coff[730 ] = 256'h00006c75ffffbc05ffffbc05ffff938bffff938b000043fb000043fb00006c75;
    assign coff[731 ] = 256'h00001c9fffff833effff833effffe361ffffe36100007cc200007cc200001c9f;
    assign coff[732 ] = 256'h000077a2ffffd27cffffd27cffff885effff885e00002d8400002d84000077a2;
    assign coff[733 ] = 256'h00003469ffff8b39ffff8b39ffffcb97ffffcb97000074c7000074c700003469;
    assign coff[734 ] = 256'h00005d1cffffa82bffffa82bffffa2e4ffffa2e4000057d5000057d500005d1c;
    assign coff[735 ] = 256'h000003bbffff800effff800efffffc45fffffc4500007ff200007ff2000003bb;
    assign coff[736 ] = 256'h00007fe0fffffa4ffffffa4fffff8020ffff8020000005b1000005b100007fe0;
    assign coff[737 ] = 256'h00005665ffffa18effffa18effffa99bffffa99b00005e7200005e7200005665;
    assign coff[738 ] = 256'h000073f6ffffc9ceffffc9ceffff8c0affff8c0a0000363200003632000073f6;
    assign coff[739 ] = 256'h00002badffff87afffff87afffffd453ffffd453000078510000785100002bad;
    assign coff[740 ] = 256'h00007c4effffe178ffffe178ffff83b2ffff83b200001e8800001e8800007c4e;
    assign coff[741 ] = 256'h0000424fffff9284ffff9284ffffbdb1ffffbdb100006d7c00006d7c0000424f;
    assign coff[742 ] = 256'h00006729ffffb439ffffb439ffff98d7ffff98d700004bc700004bc700006729;
    assign coff[743 ] = 256'h0000135dffff8179ffff8179ffffeca3ffffeca300007e8700007e870000135d;
    assign coff[744 ] = 256'h00007eb3ffffedcdffffedcdffff814dffff814d000012330000123300007eb3;
    assign coff[745 ] = 256'h00004cb9ffff998bffff998bffffb347ffffb347000066750000667500004cb9;
    assign coff[746 ] = 256'h00006e17ffffbeb3ffffbeb3ffff91e9ffff91e90000414d0000414d00006e17;
    assign coff[747 ] = 256'h00001facffff83fbffff83fbffffe054ffffe05400007c0500007c0500001fac;
    assign coff[748 ] = 256'h000078b7ffffd56fffffd56fffff8749ffff874900002a9100002a91000078b7;
    assign coff[749 ] = 256'h00003742ffff8c8bffff8c8bffffc8beffffc8be000073750000737500003742;
    assign coff[750 ] = 256'h00005f3cffffaa7affffaa7affffa0c4ffffa0c4000055860000558600005f3c;
    assign coff[751 ] = 256'h000006deffff802fffff802ffffff922fffff92200007fd100007fd1000006de;
    assign coff[752 ] = 256'h00007f71fffff40afffff40affff808fffff808f00000bf600000bf600007f71;
    assign coff[753 ] = 256'h000051a8ffff9d6effff9d6effffae58ffffae580000629200006292000051a8;
    assign coff[754 ] = 256'h0000712affffc42effffc42effff8ed6ffff8ed600003bd200003bd20000712a;
    assign coff[755 ] = 256'h000025b8ffff85afffff85afffffda48ffffda4800007a5100007a51000025b8;
    assign coff[756 ] = 256'h00007aa8ffffdb68ffffdb68ffff8558ffff8558000024980000249800007aa8;
    assign coff[757 ] = 256'h00003cdcffff8f65ffff8f65ffffc324ffffc3240000709b0000709b00003cdc;
    assign coff[758 ] = 256'h00006351ffffaf41ffffaf41ffff9cafffff9caf000050bf000050bf00006351;
    assign coff[759 ] = 256'h00000d22ffff80adffff80adfffff2defffff2de00007f5300007f5300000d22;
    assign coff[760 ] = 256'h00007da7ffffe79bffffe79bffff8259ffff8259000018650000186500007da7;
    assign coff[761 ] = 256'h0000479affff95e6ffff95e6ffffb866ffffb86600006a1a00006a1a0000479a;
    assign coff[762 ] = 256'h00006ac1ffffb961ffffb961ffff953fffff953f0000469f0000469f00006ac1;
    assign coff[763 ] = 256'h0000198dffff8293ffff8293ffffe673ffffe67300007d6d00007d6d0000198d;
    assign coff[764 ] = 256'h0000767bffffcf90ffffcf90ffff8985ffff898500003070000030700000767b;
    assign coff[765 ] = 256'h00003187ffff89f8ffff89f8ffffce79ffffce79000076080000760800003187;
    assign coff[766 ] = 256'h00005aedffffa5e8ffffa5e8ffffa513ffffa51300005a1800005a1800005aed;
    assign coff[767 ] = 256'h00000097ffff8001ffff8001ffffff69ffffff6900007fff00007fff00000097;
    assign coff[768 ] = 256'h00007fffffffff69ffffff69ffff8001ffff8001000000970000009700007fff;
    assign coff[769 ] = 256'h00005a18ffffa513ffffa513ffffa5e8ffffa5e800005aed00005aed00005a18;
    assign coff[770 ] = 256'h00007608ffffce79ffffce79ffff89f8ffff89f8000031870000318700007608;
    assign coff[771 ] = 256'h00003070ffff8985ffff8985ffffcf90ffffcf900000767b0000767b00003070;
    assign coff[772 ] = 256'h00007d6dffffe673ffffe673ffff8293ffff82930000198d0000198d00007d6d;
    assign coff[773 ] = 256'h0000469fffff953fffff953fffffb961ffffb96100006ac100006ac10000469f;
    assign coff[774 ] = 256'h00006a1affffb866ffffb866ffff95e6ffff95e60000479a0000479a00006a1a;
    assign coff[775 ] = 256'h00001865ffff8259ffff8259ffffe79bffffe79b00007da700007da700001865;
    assign coff[776 ] = 256'h00007f53fffff2defffff2deffff80adffff80ad00000d2200000d2200007f53;
    assign coff[777 ] = 256'h000050bfffff9cafffff9cafffffaf41ffffaf410000635100006351000050bf;
    assign coff[778 ] = 256'h0000709bffffc324ffffc324ffff8f65ffff8f6500003cdc00003cdc0000709b;
    assign coff[779 ] = 256'h00002498ffff8558ffff8558ffffdb68ffffdb6800007aa800007aa800002498;
    assign coff[780 ] = 256'h00007a51ffffda48ffffda48ffff85afffff85af000025b8000025b800007a51;
    assign coff[781 ] = 256'h00003bd2ffff8ed6ffff8ed6ffffc42effffc42e0000712a0000712a00003bd2;
    assign coff[782 ] = 256'h00006292ffffae58ffffae58ffff9d6effff9d6e000051a8000051a800006292;
    assign coff[783 ] = 256'h00000bf6ffff808fffff808ffffff40afffff40a00007f7100007f7100000bf6;
    assign coff[784 ] = 256'h00007fd1fffff922fffff922ffff802fffff802f000006de000006de00007fd1;
    assign coff[785 ] = 256'h00005586ffffa0c4ffffa0c4ffffaa7affffaa7a00005f3c00005f3c00005586;
    assign coff[786 ] = 256'h00007375ffffc8beffffc8beffff8c8bffff8c8b000037420000374200007375;
    assign coff[787 ] = 256'h00002a91ffff8749ffff8749ffffd56fffffd56f000078b7000078b700002a91;
    assign coff[788 ] = 256'h00007c05ffffe054ffffe054ffff83fbffff83fb00001fac00001fac00007c05;
    assign coff[789 ] = 256'h0000414dffff91e9ffff91e9ffffbeb3ffffbeb300006e1700006e170000414d;
    assign coff[790 ] = 256'h00006675ffffb347ffffb347ffff998bffff998b00004cb900004cb900006675;
    assign coff[791 ] = 256'h00001233ffff814dffff814dffffedcdffffedcd00007eb300007eb300001233;
    assign coff[792 ] = 256'h00007e87ffffeca3ffffeca3ffff8179ffff81790000135d0000135d00007e87;
    assign coff[793 ] = 256'h00004bc7ffff98d7ffff98d7ffffb439ffffb439000067290000672900004bc7;
    assign coff[794 ] = 256'h00006d7cffffbdb1ffffbdb1ffff9284ffff92840000424f0000424f00006d7c;
    assign coff[795 ] = 256'h00001e88ffff83b2ffff83b2ffffe178ffffe17800007c4e00007c4e00001e88;
    assign coff[796 ] = 256'h00007851ffffd453ffffd453ffff87afffff87af00002bad00002bad00007851;
    assign coff[797 ] = 256'h00003632ffff8c0affff8c0affffc9ceffffc9ce000073f6000073f600003632;
    assign coff[798 ] = 256'h00005e72ffffa99bffffa99bffffa18effffa18e000056650000566500005e72;
    assign coff[799 ] = 256'h000005b1ffff8020ffff8020fffffa4ffffffa4f00007fe000007fe0000005b1;
    assign coff[800 ] = 256'h00007ff2fffffc45fffffc45ffff800effff800e000003bb000003bb00007ff2;
    assign coff[801 ] = 256'h000057d5ffffa2e4ffffa2e4ffffa82bffffa82b00005d1c00005d1c000057d5;
    assign coff[802 ] = 256'h000074c7ffffcb97ffffcb97ffff8b39ffff8b390000346900003469000074c7;
    assign coff[803 ] = 256'h00002d84ffff885effff885effffd27cffffd27c000077a2000077a200002d84;
    assign coff[804 ] = 256'h00007cc2ffffe361ffffe361ffff833effff833e00001c9f00001c9f00007cc2;
    assign coff[805 ] = 256'h000043fbffff938bffff938bffffbc05ffffbc0500006c7500006c75000043fb;
    assign coff[806 ] = 256'h00006850ffffb5d1ffffb5d1ffff97b0ffff97b000004a2f00004a2f00006850;
    assign coff[807 ] = 256'h0000154dffff81c9ffff81c9ffffeab3ffffeab300007e3700007e370000154d;
    assign coff[808 ] = 256'h00007ef7ffffefbfffffefbfffff8109ffff8109000010410000104100007ef7;
    assign coff[809 ] = 256'h00004e49ffff9abbffff9abbffffb1b7ffffb1b7000065450000654500004e49;
    assign coff[810 ] = 256'h00006f14ffffc066ffffc066ffff90ecffff90ec00003f9a00003f9a00006f14;
    assign coff[811 ] = 256'h00002192ffff847bffff847bffffde6effffde6e00007b8500007b8500002192;
    assign coff[812 ] = 256'h0000795bffffd74affffd74affff86a5ffff86a5000028b6000028b60000795b;
    assign coff[813 ] = 256'h00003906ffff8d67ffff8d67ffffc6faffffc6fa000072990000729900003906;
    assign coff[814 ] = 256'h00006089ffffabf3ffffabf3ffff9f77ffff9f770000540d0000540d00006089;
    assign coff[815 ] = 256'h000008d4ffff804effff804efffff72cfffff72c00007fb200007fb2000008d4;
    assign coff[816 ] = 256'h00007f9cfffff5fffffff5ffffff8064ffff806400000a0100000a0100007f9c;
    assign coff[817 ] = 256'h00005329ffff9eb2ffff9eb2ffffacd7ffffacd70000614e0000614e00005329;
    assign coff[818 ] = 256'h00007211ffffc5edffffc5edffff8defffff8def00003a1300003a1300007211;
    assign coff[819 ] = 256'h00002797ffff8647ffff8647ffffd869ffffd869000079b9000079b900002797;
    assign coff[820 ] = 256'h00007b34ffffdd4bffffdd4bffff84ccffff84cc000022b5000022b500007b34;
    assign coff[821 ] = 256'h00003e94ffff9057ffff9057ffffc16cffffc16c00006fa900006fa900003e94;
    assign coff[822 ] = 256'h0000648bffffb0c9ffffb0c9ffff9b75ffff9b7500004f3700004f370000648b;
    assign coff[823 ] = 256'h00000f15ffff80e4ffff80e4fffff0ebfffff0eb00007f1c00007f1c00000f15;
    assign coff[824 ] = 256'h00007e03ffffe989ffffe989ffff81fdffff81fd000016770000167700007e03;
    assign coff[825 ] = 256'h00004939ffff9703ffff9703ffffb6c7ffffb6c7000068fd000068fd00004939;
    assign coff[826 ] = 256'h00006bd3ffffbb06ffffbb06ffff942dffff942d000044fa000044fa00006bd3;
    assign coff[827 ] = 256'h00001b78ffff82fbffff82fbffffe488ffffe48800007d0500007d0500001b78;
    assign coff[828 ] = 256'h00007736ffffd162ffffd162ffff88caffff88ca00002e9e00002e9e00007736;
    assign coff[829 ] = 256'h00003355ffff8abeffff8abeffffccabffffccab000075420000754200003355;
    assign coff[830 ] = 256'h00005c4cffffa750ffffa750ffffa3b4ffffa3b4000058b0000058b000005c4c;
    assign coff[831 ] = 256'h0000028dffff8007ffff8007fffffd73fffffd7300007ff900007ff90000028d;
    assign coff[832 ] = 256'h00007ffbfffffdd7fffffdd7ffff8005ffff8005000002290000022900007ffb;
    assign coff[833 ] = 256'h000058f8ffffa3faffffa3faffffa708ffffa70800005c0600005c06000058f8;
    assign coff[834 ] = 256'h0000756affffcd07ffffcd07ffff8a96ffff8a96000032f9000032f90000756a;
    assign coff[835 ] = 256'h00002efbffff88efffff88efffffd105ffffd105000077110000771100002efb;
    assign coff[836 ] = 256'h00007d1affffe4eaffffe4eaffff82e6ffff82e600001b1600001b1600007d1a;
    assign coff[837 ] = 256'h0000454fffff9463ffff9463ffffbab1ffffbab100006b9d00006b9d0000454f;
    assign coff[838 ] = 256'h00006937ffffb71affffb71affff96c9ffff96c9000048e6000048e600006937;
    assign coff[839 ] = 256'h000016daffff820effff820effffe926ffffe92600007df200007df2000016da;
    assign coff[840 ] = 256'h00007f27fffff14efffff14effff80d9ffff80d900000eb200000eb200007f27;
    assign coff[841 ] = 256'h00004f85ffff9bb3ffff9bb3ffffb07bffffb07b0000644d0000644d00004f85;
    assign coff[842 ] = 256'h00006fdaffffc1c4ffffc1c4ffff9026ffff902600003e3c00003e3c00006fda;
    assign coff[843 ] = 256'h00002316ffff84e7ffff84e7ffffdceaffffdcea00007b1900007b1900002316;
    assign coff[844 ] = 256'h000079d8ffffd8c8ffffd8c8ffff8628ffff86280000273800002738000079d8;
    assign coff[845 ] = 256'h00003a6dffff8e1dffff8e1dffffc593ffffc593000071e3000071e300003a6d;
    assign coff[846 ] = 256'h00006190ffffad24ffffad24ffff9e70ffff9e70000052dc000052dc00006190;
    assign coff[847 ] = 256'h00000a65ffff806cffff806cfffff59bfffff59b00007f9400007f9400000a65;
    assign coff[848 ] = 256'h00007fb9fffff790fffff790ffff8047ffff8047000008700000087000007fb9;
    assign coff[849 ] = 256'h00005459ffff9fb9ffff9fb9ffffaba7ffffaba7000060470000604700005459;
    assign coff[850 ] = 256'h000072c5ffffc754ffffc754ffff8d3bffff8d3b000038ac000038ac000072c5;
    assign coff[851 ] = 256'h00002915ffff86c6ffff86c6ffffd6ebffffd6eb0000793a0000793a00002915;
    assign coff[852 ] = 256'h00007b9fffffdecfffffdecfffff8461ffff8461000021310000213100007b9f;
    assign coff[853 ] = 256'h00003ff1ffff911effff911effffc00fffffc00f00006ee200006ee200003ff1;
    assign coff[854 ] = 256'h00006582ffffb207ffffb207ffff9a7effff9a7e00004df900004df900006582;
    assign coff[855 ] = 256'h000010a4ffff8116ffff8116ffffef5cffffef5c00007eea00007eea000010a4;
    assign coff[856 ] = 256'h00007e48ffffeb16ffffeb16ffff81b8ffff81b8000014ea000014ea00007e48;
    assign coff[857 ] = 256'h00004a81ffff97ebffff97ebffffb57fffffb57f000068150000681500004a81;
    assign coff[858 ] = 256'h00006caaffffbc5affffbc5affff9356ffff9356000043a6000043a600006caa;
    assign coff[859 ] = 256'h00001d01ffff8354ffff8354ffffe2ffffffe2ff00007cac00007cac00001d01;
    assign coff[860 ] = 256'h000077c6ffffd2daffffd2daffff883affff883a00002d2600002d26000077c6;
    assign coff[861 ] = 256'h000034c4ffff8b62ffff8b62ffffcb3cffffcb3c0000749e0000749e000034c4;
    assign coff[862 ] = 256'h00005d61ffffa874ffffa874ffffa29fffffa29f0000578c0000578c00005d61;
    assign coff[863 ] = 256'h0000041fffff8011ffff8011fffffbe1fffffbe100007fef00007fef0000041f;
    assign coff[864 ] = 256'h00007fe4fffffab3fffffab3ffff801cffff801c0000054d0000054d00007fe4;
    assign coff[865 ] = 256'h000056afffffa1d2ffffa1d2ffffa951ffffa95100005e2e00005e2e000056af;
    assign coff[866 ] = 256'h00007421ffffca29ffffca29ffff8bdfffff8bdf000035d7000035d700007421;
    assign coff[867 ] = 256'h00002c0cffff87d1ffff87d1ffffd3f4ffffd3f40000782f0000782f00002c0c;
    assign coff[868 ] = 256'h00007c66ffffe1daffffe1daffff839affff839a00001e2600001e2600007c66;
    assign coff[869 ] = 256'h000042a5ffff92b8ffff92b8ffffbd5bffffbd5b00006d4800006d48000042a5;
    assign coff[870 ] = 256'h00006764ffffb48bffffb48bffff989cffff989c00004b7500004b7500006764;
    assign coff[871 ] = 256'h000013c1ffff8188ffff8188ffffec3fffffec3f00007e7800007e78000013c1;
    assign coff[872 ] = 256'h00007ec1ffffee31ffffee31ffff813fffff813f000011cf000011cf00007ec1;
    assign coff[873 ] = 256'h00004d09ffff99c7ffff99c7ffffb2f7ffffb2f7000066390000663900004d09;
    assign coff[874 ] = 256'h00006e4affffbf0affffbf0affff91b6ffff91b6000040f6000040f600006e4a;
    assign coff[875 ] = 256'h0000200effff8414ffff8414ffffdff2ffffdff200007bec00007bec0000200e;
    assign coff[876 ] = 256'h000078d8ffffd5ceffffd5ceffff8728ffff872800002a3200002a32000078d8;
    assign coff[877 ] = 256'h0000379dffff8cb6ffff8cb6ffffc863ffffc8630000734a0000734a0000379d;
    assign coff[878 ] = 256'h00005f80ffffaac5ffffaac5ffffa080ffffa0800000553b0000553b00005f80;
    assign coff[879 ] = 256'h00000743ffff8035ffff8035fffff8bdfffff8bd00007fcb00007fcb00000743;
    assign coff[880 ] = 256'h00007f7afffff46efffff46effff8086ffff808600000b9200000b9200007f7a;
    assign coff[881 ] = 256'h000051f5ffff9daeffff9daeffffae0bffffae0b0000625200006252000051f5;
    assign coff[882 ] = 256'h00007158ffffc487ffffc487ffff8ea8ffff8ea800003b7900003b7900007158;
    assign coff[883 ] = 256'h00002618ffff85cdffff85cdffffd9e8ffffd9e800007a3300007a3300002618;
    assign coff[884 ] = 256'h00007ac5ffffdbc9ffffdbc9ffff853bffff853b000024370000243700007ac5;
    assign coff[885 ] = 256'h00003d34ffff8f95ffff8f95ffffc2ccffffc2cc0000706b0000706b00003d34;
    assign coff[886 ] = 256'h00006391ffffaf8fffffaf8fffff9c6fffff9c6f000050710000507100006391;
    assign coff[887 ] = 256'h00000d86ffff80b7ffff80b7fffff27afffff27a00007f4900007f4900000d86;
    assign coff[888 ] = 256'h00007dbaffffe7feffffe7feffff8246ffff8246000018020000180200007dba;
    assign coff[889 ] = 256'h000047edffff961fffff961fffffb813ffffb813000069e1000069e1000047ed;
    assign coff[890 ] = 256'h00006af8ffffb9b5ffffb9b5ffff9508ffff95080000464b0000464b00006af8;
    assign coff[891 ] = 256'h000019efffff82a8ffff82a8ffffe611ffffe61100007d5800007d58000019ef;
    assign coff[892 ] = 256'h000076a1ffffcfedffffcfedffff895fffff895f0000301300003013000076a1;
    assign coff[893 ] = 256'h000031e4ffff8a1fffff8a1fffffce1cffffce1c000075e1000075e1000031e4;
    assign coff[894 ] = 256'h00005b34ffffa630ffffa630ffffa4ccffffa4cc000059d0000059d000005b34;
    assign coff[895 ] = 256'h000000fbffff8001ffff8001ffffff05ffffff0500007fff00007fff000000fb;
    assign coff[896 ] = 256'h00007ffefffffea0fffffea0ffff8002ffff8002000001600000016000007ffe;
    assign coff[897 ] = 256'h00005988ffffa486ffffa486ffffa678ffffa67800005b7a00005b7a00005988;
    assign coff[898 ] = 256'h000075b9ffffcdc0ffffcdc0ffff8a47ffff8a470000324000003240000075b9;
    assign coff[899 ] = 256'h00002fb6ffff8939ffff8939ffffd04affffd04a000076c7000076c700002fb6;
    assign coff[900 ] = 256'h00007d44ffffe5afffffe5afffff82bcffff82bc00001a5100001a5100007d44;
    assign coff[901 ] = 256'h000045f7ffff94d0ffff94d0ffffba09ffffba0900006b3000006b30000045f7;
    assign coff[902 ] = 256'h000069a9ffffb7c0ffffb7c0ffff9657ffff96570000484000004840000069a9;
    assign coff[903 ] = 256'h0000179fffff8233ffff8233ffffe861ffffe86100007dcd00007dcd0000179f;
    assign coff[904 ] = 256'h00007f3efffff216fffff216ffff80c2ffff80c200000dea00000dea00007f3e;
    assign coff[905 ] = 256'h00005023ffff9c30ffff9c30ffffafddffffafdd000063d0000063d000005023;
    assign coff[906 ] = 256'h0000703bffffc274ffffc274ffff8fc5ffff8fc500003d8c00003d8c0000703b;
    assign coff[907 ] = 256'h000023d7ffff851fffff851fffffdc29ffffdc2900007ae100007ae1000023d7;
    assign coff[908 ] = 256'h00007a15ffffd988ffffd988ffff85ebffff85eb000026780000267800007a15;
    assign coff[909 ] = 256'h00003b20ffff8e79ffff8e79ffffc4e0ffffc4e0000071870000718700003b20;
    assign coff[910 ] = 256'h00006211ffffadbdffffadbdffff9defffff9def000052430000524300006211;
    assign coff[911 ] = 256'h00000b2dffff807dffff807dfffff4d3fffff4d300007f8300007f8300000b2d;
    assign coff[912 ] = 256'h00007fc5fffff859fffff859ffff803bffff803b000007a7000007a700007fc5;
    assign coff[913 ] = 256'h000054f0ffffa03effffa03effffab10ffffab1000005fc200005fc2000054f0;
    assign coff[914 ] = 256'h0000731effffc809ffffc809ffff8ce2ffff8ce2000037f7000037f70000731e;
    assign coff[915 ] = 256'h000029d3ffff8707ffff8707ffffd62dffffd62d000078f9000078f9000029d3;
    assign coff[916 ] = 256'h00007bd3ffffdf91ffffdf91ffff842dffff842d0000206f0000206f00007bd3;
    assign coff[917 ] = 256'h0000409fffff9183ffff9183ffffbf61ffffbf6100006e7d00006e7d0000409f;
    assign coff[918 ] = 256'h000065fcffffb2a7ffffb2a7ffff9a04ffff9a0400004d5900004d59000065fc;
    assign coff[919 ] = 256'h0000116cffff8131ffff8131ffffee94ffffee9400007ecf00007ecf0000116c;
    assign coff[920 ] = 256'h00007e68ffffebdcffffebdcffff8198ffff8198000014240000142400007e68;
    assign coff[921 ] = 256'h00004b24ffff9860ffff9860ffffb4dcffffb4dc000067a0000067a000004b24;
    assign coff[922 ] = 256'h00006d14ffffbd05ffffbd05ffff92ecffff92ec000042fb000042fb00006d14;
    assign coff[923 ] = 256'h00001dc4ffff8382ffff8382ffffe23cffffe23c00007c7e00007c7e00001dc4;
    assign coff[924 ] = 256'h0000780cffffd396ffffd396ffff87f4ffff87f400002c6a00002c6a0000780c;
    assign coff[925 ] = 256'h0000357bffff8bb5ffff8bb5ffffca85ffffca850000744b0000744b0000357b;
    assign coff[926 ] = 256'h00005deaffffa907ffffa907ffffa216ffffa216000056f9000056f900005dea;
    assign coff[927 ] = 256'h000004e8ffff8018ffff8018fffffb18fffffb1800007fe800007fe8000004e8;
    assign coff[928 ] = 256'h00007fecfffffb7cfffffb7cffff8014ffff8014000004840000048400007fec;
    assign coff[929 ] = 256'h00005743ffffa25bffffa25bffffa8bdffffa8bd00005da500005da500005743;
    assign coff[930 ] = 256'h00007475ffffcae0ffffcae0ffff8b8bffff8b8b000035200000352000007475;
    assign coff[931 ] = 256'h00002cc8ffff8817ffff8817ffffd338ffffd338000077e9000077e900002cc8;
    assign coff[932 ] = 256'h00007c95ffffe29effffe29effff836bffff836b00001d6200001d6200007c95;
    assign coff[933 ] = 256'h00004351ffff9321ffff9321ffffbcafffffbcaf00006cdf00006cdf00004351;
    assign coff[934 ] = 256'h000067daffffb52dffffb52dffff9826ffff982600004ad300004ad3000067da;
    assign coff[935 ] = 256'h00001487ffff81a8ffff81a8ffffeb79ffffeb7900007e5800007e5800001487;
    assign coff[936 ] = 256'h00007eddffffeef8ffffeef8ffff8123ffff8123000011080000110800007edd;
    assign coff[937 ] = 256'h00004da9ffff9a40ffff9a40ffffb257ffffb257000065c0000065c000004da9;
    assign coff[938 ] = 256'h00006eb0ffffbfb8ffffbfb8ffff9150ffff9150000040480000404800006eb0;
    assign coff[939 ] = 256'h000020d0ffff8447ffff8447ffffdf30ffffdf3000007bb900007bb9000020d0;
    assign coff[940 ] = 256'h0000791affffd68cffffd68cffff86e6ffff86e600002974000029740000791a;
    assign coff[941 ] = 256'h00003852ffff8d0effff8d0effffc7aeffffc7ae000072f2000072f200003852;
    assign coff[942 ] = 256'h00006005ffffab5cffffab5cffff9ffbffff9ffb000054a4000054a400006005;
    assign coff[943 ] = 256'h0000080cffff8041ffff8041fffff7f4fffff7f400007fbf00007fbf0000080c;
    assign coff[944 ] = 256'h00007f8bfffff537fffff537ffff8075ffff807500000ac900000ac900007f8b;
    assign coff[945 ] = 256'h00005290ffff9e2fffff9e2fffffad70ffffad70000061d1000061d100005290;
    assign coff[946 ] = 256'h000071b5ffffc53affffc53affff8e4bffff8e4b00003ac600003ac6000071b5;
    assign coff[947 ] = 256'h000026d8ffff8609ffff8609ffffd928ffffd928000079f7000079f7000026d8;
    assign coff[948 ] = 256'h00007afdffffdc8affffdc8affff8503ffff8503000023760000237600007afd;
    assign coff[949 ] = 256'h00003de4ffff8ff5ffff8ff5ffffc21cffffc21c0000700b0000700b00003de4;
    assign coff[950 ] = 256'h0000640fffffb02cffffb02cffff9bf1ffff9bf100004fd400004fd40000640f;
    assign coff[951 ] = 256'h00000e4effff80cdffff80cdfffff1b2fffff1b200007f3300007f3300000e4e;
    assign coff[952 ] = 256'h00007de0ffffe8c4ffffe8c4ffff8220ffff82200000173c0000173c00007de0;
    assign coff[953 ] = 256'h00004893ffff9690ffff9690ffffb76dffffb76d000069700000697000004893;
    assign coff[954 ] = 256'h00006b66ffffba5dffffba5dffff949affff949a000045a3000045a300006b66;
    assign coff[955 ] = 256'h00001ab4ffff82d1ffff82d1ffffe54cffffe54c00007d2f00007d2f00001ab4;
    assign coff[956 ] = 256'h000076ecffffd0a7ffffd0a7ffff8914ffff891400002f5900002f59000076ec;
    assign coff[957 ] = 256'h0000329dffff8a6effff8a6effffcd63ffffcd6300007592000075920000329d;
    assign coff[958 ] = 256'h00005bc0ffffa6c0ffffa6c0ffffa440ffffa440000059400000594000005bc0;
    assign coff[959 ] = 256'h000001c4ffff8003ffff8003fffffe3cfffffe3c00007ffd00007ffd000001c4;
    assign coff[960 ] = 256'h00007ff7fffffd0efffffd0effff8009ffff8009000002f2000002f200007ff7;
    assign coff[961 ] = 256'h00005867ffffa36fffffa36fffffa799ffffa79900005c9100005c9100005867;
    assign coff[962 ] = 256'h00007519ffffcc4fffffcc4fffff8ae7ffff8ae7000033b1000033b100007519;
    assign coff[963 ] = 256'h00002e40ffff88a6ffff88a6ffffd1c0ffffd1c00000775a0000775a00002e40;
    assign coff[964 ] = 256'h00007cefffffe426ffffe426ffff8311ffff831100001bda00001bda00007cef;
    assign coff[965 ] = 256'h000044a5ffff93f7ffff93f7ffffbb5bffffbb5b00006c0900006c09000044a5;
    assign coff[966 ] = 256'h000068c4ffffb675ffffb675ffff973cffff973c0000498b0000498b000068c4;
    assign coff[967 ] = 256'h00001614ffff81ebffff81ebffffe9ecffffe9ec00007e1500007e1500001614;
    assign coff[968 ] = 256'h00007f10fffff087fffff087ffff80f0ffff80f000000f7900000f7900007f10;
    assign coff[969 ] = 256'h00004ee8ffff9b36ffff9b36ffffb118ffffb118000064ca000064ca00004ee8;
    assign coff[970 ] = 256'h00006f78ffffc114ffffc114ffff9088ffff908800003eec00003eec00006f78;
    assign coff[971 ] = 256'h00002254ffff84b0ffff84b0ffffddacffffddac00007b5000007b5000002254;
    assign coff[972 ] = 256'h0000799affffd809ffffd809ffff8666ffff8666000027f7000027f70000799a;
    assign coff[973 ] = 256'h000039baffff8dc1ffff8dc1ffffc646ffffc6460000723f0000723f000039ba;
    assign coff[974 ] = 256'h0000610dffffac8bffffac8bffff9ef3ffff9ef300005375000053750000610d;
    assign coff[975 ] = 256'h0000099dffff805dffff805dfffff663fffff66300007fa300007fa30000099d;
    assign coff[976 ] = 256'h00007fabfffff6c8fffff6c8ffff8055ffff8055000009380000093800007fab;
    assign coff[977 ] = 256'h000053c1ffff9f35ffff9f35ffffac3fffffac3f000060cb000060cb000053c1;
    assign coff[978 ] = 256'h0000726cffffc6a0ffffc6a0ffff8d94ffff8d9400003960000039600000726c;
    assign coff[979 ] = 256'h00002856ffff8686ffff8686ffffd7aaffffd7aa0000797a0000797a00002856;
    assign coff[980 ] = 256'h00007b6affffde0dffffde0dffff8496ffff8496000021f3000021f300007b6a;
    assign coff[981 ] = 256'h00003f43ffff90baffff90baffffc0bdffffc0bd00006f4600006f4600003f43;
    assign coff[982 ] = 256'h00006507ffffb168ffffb168ffff9af9ffff9af900004e9800004e9800006507;
    assign coff[983 ] = 256'h00000fddffff80fdffff80fdfffff023fffff02300007f0300007f0300000fdd;
    assign coff[984 ] = 256'h00007e26ffffea4fffffea4fffff81daffff81da000015b1000015b100007e26;
    assign coff[985 ] = 256'h000049ddffff9776ffff9776ffffb623ffffb6230000688a0000688a000049dd;
    assign coff[986 ] = 256'h00006c3fffffbbb0ffffbbb0ffff93c1ffff93c1000044500000445000006c3f;
    assign coff[987 ] = 256'h00001c3dffff8327ffff8327ffffe3c3ffffe3c300007cd900007cd900001c3d;
    assign coff[988 ] = 256'h0000777effffd21effffd21effff8882ffff888200002de200002de20000777e;
    assign coff[989 ] = 256'h0000340dffff8b10ffff8b10ffffcbf3ffffcbf3000074f0000074f00000340d;
    assign coff[990 ] = 256'h00005cd7ffffa7e2ffffa7e2ffffa329ffffa3290000581e0000581e00005cd7;
    assign coff[991 ] = 256'h00000356ffff800bffff800bfffffcaafffffcaa00007ff500007ff500000356;
    assign coff[992 ] = 256'h00007fdbfffff9eafffff9eaffff8025ffff8025000006160000061600007fdb;
    assign coff[993 ] = 256'h0000561bffffa14affffa14affffa9e5ffffa9e500005eb600005eb60000561b;
    assign coff[994 ] = 256'h000073cbffffc973ffffc973ffff8c35ffff8c350000368d0000368d000073cb;
    assign coff[995 ] = 256'h00002b4fffff878cffff878cffffd4b1ffffd4b1000078740000787400002b4f;
    assign coff[996 ] = 256'h00007c36ffffe117ffffe117ffff83caffff83ca00001ee900001ee900007c36;
    assign coff[997 ] = 256'h000041f9ffff9250ffff9250ffffbe07ffffbe0700006db000006db0000041f9;
    assign coff[998 ] = 256'h000066edffffb3e9ffffb3e9ffff9913ffff991300004c1700004c17000066ed;
    assign coff[999 ] = 256'h000012faffff816affff816affffed06ffffed0600007e9600007e96000012fa;
    assign coff[1000] = 256'h00007ea5ffffed6affffed6affff815bffff815b000012960000129600007ea5;
    assign coff[1001] = 256'h00004c68ffff994effff994effffb398ffffb398000066b2000066b200004c68;
    assign coff[1002] = 256'h00006de4ffffbe5dffffbe5dffff921cffff921c000041a3000041a300006de4;
    assign coff[1003] = 256'h00001f4bffff83e2ffff83e2ffffe0b5ffffe0b500007c1e00007c1e00001f4b;
    assign coff[1004] = 256'h00007895ffffd510ffffd510ffff876bffff876b00002af000002af000007895;
    assign coff[1005] = 256'h000036e8ffff8c60ffff8c60ffffc918ffffc918000073a0000073a0000036e8;
    assign coff[1006] = 256'h00005ef9ffffaa30ffffaa30ffffa107ffffa107000055d0000055d000005ef9;
    assign coff[1007] = 256'h0000067affff802affff802afffff986fffff98600007fd600007fd60000067a;
    assign coff[1008] = 256'h00007f67fffff3a6fffff3a6ffff8099ffff809900000c5a00000c5a00007f67;
    assign coff[1009] = 256'h0000515bffff9d2effff9d2effffaea5ffffaea5000062d2000062d20000515b;
    assign coff[1010] = 256'h000070faffffc3d6ffffc3d6ffff8f06ffff8f0600003c2a00003c2a000070fa;
    assign coff[1011] = 256'h00002558ffff8592ffff8592ffffdaa8ffffdaa800007a6e00007a6e00002558;
    assign coff[1012] = 256'h00007a8cffffdb08ffffdb08ffff8574ffff8574000024f8000024f800007a8c;
    assign coff[1013] = 256'h00003c83ffff8f35ffff8f35ffffc37dffffc37d000070cb000070cb00003c83;
    assign coff[1014] = 256'h00006312ffffaef3ffffaef3ffff9ceeffff9cee0000510d0000510d00006312;
    assign coff[1015] = 256'h00000cbeffff80a3ffff80a3fffff342fffff34200007f5d00007f5d00000cbe;
    assign coff[1016] = 256'h00007d94ffffe739ffffe739ffff826cffff826c000018c7000018c700007d94;
    assign coff[1017] = 256'h00004747ffff95aeffff95aeffffb8b9ffffb8b900006a5200006a5200004747;
    assign coff[1018] = 256'h00006a89ffffb90dffffb90dffff9577ffff9577000046f3000046f300006a89;
    assign coff[1019] = 256'h0000192affff827fffff827fffffe6d6ffffe6d600007d8100007d810000192a;
    assign coff[1020] = 256'h00007655ffffcf33ffffcf33ffff89abffff89ab000030cd000030cd00007655;
    assign coff[1021] = 256'h0000312affff89d2ffff89d2ffffced6ffffced60000762e0000762e0000312a;
    assign coff[1022] = 256'h00005aa6ffffa5a1ffffa5a1ffffa55affffa55a00005a5f00005a5f00005aa6;
    assign coff[1023] = 256'h00000032ffff8001ffff8001ffffffceffffffce00007fff00007fff00000032;
    assign coff[1024] = 256'h00007fffffffffe7ffffffe7ffff8001ffff8001000000190000001900007fff;
    assign coff[1025] = 256'h00005a71ffffa56cffffa56cffffa58fffffa58f00005a9400005a9400005a71;
    assign coff[1026] = 256'h00007638ffffceedffffceedffff89c8ffff89c8000031130000311300007638;
    assign coff[1027] = 256'h000030e5ffff89b5ffff89b5ffffcf1bffffcf1b0000764b0000764b000030e5;
    assign coff[1028] = 256'h00007d85ffffe6efffffe6efffff827bffff827b000019110000191100007d85;
    assign coff[1029] = 256'h00004708ffff9584ffff9584ffffb8f8ffffb8f800006a7c00006a7c00004708;
    assign coff[1030] = 256'h00006a60ffffb8ceffffb8ceffff95a0ffff95a0000047320000473200006a60;
    assign coff[1031] = 256'h000018e0ffff8271ffff8271ffffe720ffffe72000007d8f00007d8f000018e0;
    assign coff[1032] = 256'h00007f60fffff35bfffff35bffff80a0ffff80a000000ca500000ca500007f60;
    assign coff[1033] = 256'h00005120ffff9cfeffff9cfeffffaee0ffffaee0000063020000630200005120;
    assign coff[1034] = 256'h000070d7ffffc393ffffc393ffff8f29ffff8f2900003c6d00003c6d000070d7;
    assign coff[1035] = 256'h00002510ffff857cffff857cffffdaf0ffffdaf000007a8400007a8400002510;
    assign coff[1036] = 256'h00007a76ffffdac0ffffdac0ffff858affff858a000025400000254000007a76;
    assign coff[1037] = 256'h00003c41ffff8f11ffff8f11ffffc3bfffffc3bf000070ef000070ef00003c41;
    assign coff[1038] = 256'h000062e2ffffaeb9ffffaeb9ffff9d1effff9d1e0000514700005147000062e2;
    assign coff[1039] = 256'h00000c73ffff809bffff809bfffff38dfffff38d00007f6500007f6500000c73;
    assign coff[1040] = 256'h00007fd7fffff99ffffff99fffff8029ffff8029000006610000066100007fd7;
    assign coff[1041] = 256'h000055e3ffffa118ffffa118ffffaa1dffffaa1d00005ee800005ee8000055e3;
    assign coff[1042] = 256'h000073abffffc92fffffc92fffff8c55ffff8c55000036d1000036d1000073ab;
    assign coff[1043] = 256'h00002b08ffff8773ffff8773ffffd4f8ffffd4f80000788d0000788d00002b08;
    assign coff[1044] = 256'h00007c24ffffe0ceffffe0ceffff83dcffff83dc00001f3200001f3200007c24;
    assign coff[1045] = 256'h000041b9ffff9229ffff9229ffffbe47ffffbe4700006dd700006dd7000041b9;
    assign coff[1046] = 256'h000066c1ffffb3acffffb3acffff993fffff993f00004c5400004c54000066c1;
    assign coff[1047] = 256'h000012afffff815fffff815fffffed51ffffed5100007ea100007ea1000012af;
    assign coff[1048] = 256'h00007e9affffed1fffffed1fffff8166ffff8166000012e1000012e100007e9a;
    assign coff[1049] = 256'h00004c2cffff9922ffff9922ffffb3d4ffffb3d4000066de000066de00004c2c;
    assign coff[1050] = 256'h00006dbdffffbe1cffffbe1cffff9243ffff9243000041e4000041e400006dbd;
    assign coff[1051] = 256'h00001f02ffff83d0ffff83d0ffffe0feffffe0fe00007c3000007c3000001f02;
    assign coff[1052] = 256'h0000787cffffd4c9ffffd4c9ffff8784ffff878400002b3700002b370000787c;
    assign coff[1053] = 256'h000036a3ffff8c3fffff8c3fffffc95dffffc95d000073c1000073c1000036a3;
    assign coff[1054] = 256'h00005ec7ffffa9f8ffffa9f8ffffa139ffffa139000056080000560800005ec7;
    assign coff[1055] = 256'h0000062fffff8026ffff8026fffff9d1fffff9d100007fda00007fda0000062f;
    assign coff[1056] = 256'h00007ff6fffffcc3fffffcc3ffff800affff800a0000033d0000033d00007ff6;
    assign coff[1057] = 256'h00005831ffffa33bffffa33bffffa7cfffffa7cf00005cc500005cc500005831;
    assign coff[1058] = 256'h000074fbffffcc0affffcc0affff8b05ffff8b05000033f6000033f6000074fb;
    assign coff[1059] = 256'h00002dfaffff888bffff888bffffd206ffffd206000077750000777500002dfa;
    assign coff[1060] = 256'h00007cdeffffe3dcffffe3dcffff8322ffff832200001c2400001c2400007cde;
    assign coff[1061] = 256'h00004466ffff93ceffff93ceffffbb9affffbb9a00006c3200006c3200004466;
    assign coff[1062] = 256'h00006898ffffb637ffffb637ffff9768ffff9768000049c9000049c900006898;
    assign coff[1063] = 256'h000015c9ffff81deffff81deffffea37ffffea3700007e2200007e22000015c9;
    assign coff[1064] = 256'h00007f06fffff03cfffff03cffff80faffff80fa00000fc400000fc400007f06;
    assign coff[1065] = 256'h00004eacffff9b08ffff9b08ffffb154ffffb154000064f8000064f800004eac;
    assign coff[1066] = 256'h00006f53ffffc0d3ffffc0d3ffff90adffff90ad00003f2d00003f2d00006f53;
    assign coff[1067] = 256'h0000220bffff849cffff849cffffddf5ffffddf500007b6400007b640000220b;
    assign coff[1068] = 256'h00007982ffffd7c1ffffd7c1ffff867effff867e0000283f0000283f00007982;
    assign coff[1069] = 256'h00003976ffff8da0ffff8da0ffffc68affffc68a000072600000726000003976;
    assign coff[1070] = 256'h000060dcffffac52ffffac52ffff9f24ffff9f24000053ae000053ae000060dc;
    assign coff[1071] = 256'h00000951ffff8057ffff8057fffff6affffff6af00007fa900007fa900000951;
    assign coff[1072] = 256'h00007fa5fffff67cfffff67cffff805bffff805b000009840000098400007fa5;
    assign coff[1073] = 256'h00005388ffff9f03ffff9f03ffffac78ffffac78000060fd000060fd00005388;
    assign coff[1074] = 256'h0000724affffc65dffffc65dffff8db6ffff8db6000039a3000039a30000724a;
    assign coff[1075] = 256'h0000280fffff866effff866effffd7f1ffffd7f100007992000079920000280f;
    assign coff[1076] = 256'h00007b56ffffddc4ffffddc4ffff84aaffff84aa0000223c0000223c00007b56;
    assign coff[1077] = 256'h00003f01ffff9095ffff9095ffffc0ffffffc0ff00006f6b00006f6b00003f01;
    assign coff[1078] = 256'h000064d9ffffb12cffffb12cffff9b27ffff9b2700004ed400004ed4000064d9;
    assign coff[1079] = 256'h00000f92ffff80f3ffff80f3fffff06efffff06e00007f0d00007f0d00000f92;
    assign coff[1080] = 256'h00007e19ffffea05ffffea05ffff81e7ffff81e7000015fb000015fb00007e19;
    assign coff[1081] = 256'h000049a0ffff974bffff974bffffb660ffffb660000068b5000068b5000049a0;
    assign coff[1082] = 256'h00006c17ffffbb70ffffbb70ffff93e9ffff93e9000044900000449000006c17;
    assign coff[1083] = 256'h00001bf3ffff8317ffff8317ffffe40dffffe40d00007ce900007ce900001bf3;
    assign coff[1084] = 256'h00007763ffffd1d8ffffd1d8ffff889dffff889d00002e2800002e2800007763;
    assign coff[1085] = 256'h000033c8ffff8af1ffff8af1ffffcc38ffffcc380000750f0000750f000033c8;
    assign coff[1086] = 256'h00005ca3ffffa7abffffa7abffffa35dffffa35d000058550000585500005ca3;
    assign coff[1087] = 256'h0000030bffff8009ffff8009fffffcf5fffffcf500007ff700007ff70000030b;
    assign coff[1088] = 256'h00007ffdfffffe55fffffe55ffff8003ffff8003000001ab000001ab00007ffd;
    assign coff[1089] = 256'h00005952ffffa451ffffa451ffffa6aeffffa6ae00005baf00005baf00005952;
    assign coff[1090] = 256'h0000759cffffcd7bffffcd7bffff8a64ffff8a6400003285000032850000759c;
    assign coff[1091] = 256'h00002f70ffff891dffff891dffffd090ffffd090000076e3000076e300002f70;
    assign coff[1092] = 256'h00007d34ffffe565ffffe565ffff82ccffff82cc00001a9b00001a9b00007d34;
    assign coff[1093] = 256'h000045b8ffff94a7ffff94a7ffffba48ffffba4800006b5900006b59000045b8;
    assign coff[1094] = 256'h0000697effffb781ffffb781ffff9682ffff96820000487f0000487f0000697e;
    assign coff[1095] = 256'h00001755ffff8225ffff8225ffffe8abffffe8ab00007ddb00007ddb00001755;
    assign coff[1096] = 256'h00007f36fffff1cbfffff1cbffff80caffff80ca00000e3500000e3500007f36;
    assign coff[1097] = 256'h00004fe8ffff9c01ffff9c01ffffb018ffffb018000063ff000063ff00004fe8;
    assign coff[1098] = 256'h00007017ffffc232ffffc232ffff8fe9ffff8fe900003dce00003dce00007017;
    assign coff[1099] = 256'h0000238effff850affff850affffdc72ffffdc7200007af600007af60000238e;
    assign coff[1100] = 256'h000079feffffd940ffffd940ffff8602ffff8602000026c0000026c0000079fe;
    assign coff[1101] = 256'h00003addffff8e56ffff8e56ffffc523ffffc523000071aa000071aa00003add;
    assign coff[1102] = 256'h000061e1ffffad84ffffad84ffff9e1fffff9e1f0000527c0000527c000061e1;
    assign coff[1103] = 256'h00000ae2ffff8077ffff8077fffff51efffff51e00007f8900007f8900000ae2;
    assign coff[1104] = 256'h00007fc1fffff80efffff80effff803fffff803f000007f2000007f200007fc1;
    assign coff[1105] = 256'h000054b7ffffa00cffffa00cffffab49ffffab4900005ff400005ff4000054b7;
    assign coff[1106] = 256'h000072fdffffc7c5ffffc7c5ffff8d03ffff8d030000383b0000383b000072fd;
    assign coff[1107] = 256'h0000298cffff86eeffff86eeffffd674ffffd67400007912000079120000298c;
    assign coff[1108] = 256'h00007bbfffffdf48ffffdf48ffff8441ffff8441000020b8000020b800007bbf;
    assign coff[1109] = 256'h0000405effff915dffff915dffffbfa2ffffbfa200006ea300006ea30000405e;
    assign coff[1110] = 256'h000065cfffffb26bffffb26bffff9a31ffff9a3100004d9500004d95000065cf;
    assign coff[1111] = 256'h00001121ffff8127ffff8127ffffeedfffffeedf00007ed900007ed900001121;
    assign coff[1112] = 256'h00007e5cffffeb92ffffeb92ffff81a4ffff81a40000146e0000146e00007e5c;
    assign coff[1113] = 256'h00004ae7ffff9834ffff9834ffffb519ffffb519000067cc000067cc00004ae7;
    assign coff[1114] = 256'h00006cecffffbcc5ffffbcc5ffff9314ffff93140000433b0000433b00006cec;
    assign coff[1115] = 256'h00001d7bffff8371ffff8371ffffe285ffffe28500007c8f00007c8f00001d7b;
    assign coff[1116] = 256'h000077f2ffffd34fffffd34fffff880effff880e00002cb100002cb1000077f2;
    assign coff[1117] = 256'h00003537ffff8b96ffff8b96ffffcac9ffffcac90000746a0000746a00003537;
    assign coff[1118] = 256'h00005db7ffffa8d0ffffa8d0ffffa249ffffa249000057300000573000005db7;
    assign coff[1119] = 256'h0000049dffff8015ffff8015fffffb63fffffb6300007feb00007feb0000049d;
    assign coff[1120] = 256'h00007fe9fffffb31fffffb31ffff8017ffff8017000004cf000004cf00007fe9;
    assign coff[1121] = 256'h0000570cffffa227ffffa227ffffa8f4ffffa8f400005dd900005dd90000570c;
    assign coff[1122] = 256'h00007455ffffca9cffffca9cffff8babffff8bab000035640000356400007455;
    assign coff[1123] = 256'h00002c81ffff87fdffff87fdffffd37fffffd37f000078030000780300002c81;
    assign coff[1124] = 256'h00007c83ffffe254ffffe254ffff837dffff837d00001dac00001dac00007c83;
    assign coff[1125] = 256'h00004310ffff92faffff92faffffbcf0ffffbcf000006d0600006d0600004310;
    assign coff[1126] = 256'h000067aeffffb4f0ffffb4f0ffff9852ffff985200004b1000004b10000067ae;
    assign coff[1127] = 256'h0000143dffff819cffff819cffffebc3ffffebc300007e6400007e640000143d;
    assign coff[1128] = 256'h00007ed3ffffeeadffffeeadffff812dffff812d000011530000115300007ed3;
    assign coff[1129] = 256'h00004d6dffff9a13ffff9a13ffffb293ffffb293000065ed000065ed00004d6d;
    assign coff[1130] = 256'h00006e8affffbf76ffffbf76ffff9176ffff91760000408a0000408a00006e8a;
    assign coff[1131] = 256'h00002087ffff8434ffff8434ffffdf79ffffdf7900007bcc00007bcc00002087;
    assign coff[1132] = 256'h00007901ffffd644ffffd644ffff86ffffff86ff000029bc000029bc00007901;
    assign coff[1133] = 256'h0000380effff8cedffff8cedffffc7f2ffffc7f200007313000073130000380e;
    assign coff[1134] = 256'h00005fd3ffffab23ffffab23ffffa02dffffa02d000054dd000054dd00005fd3;
    assign coff[1135] = 256'h000007c0ffff803cffff803cfffff840fffff84000007fc400007fc4000007c0;
    assign coff[1136] = 256'h00007f85fffff4ecfffff4ecffff807bffff807b00000b1400000b1400007f85;
    assign coff[1137] = 256'h00005256ffff9dffffff9dffffffadaaffffadaa000062010000620100005256;
    assign coff[1138] = 256'h00007193ffffc4f7ffffc4f7ffff8e6dffff8e6d00003b0900003b0900007193;
    assign coff[1139] = 256'h00002690ffff85f2ffff85f2ffffd970ffffd97000007a0e00007a0e00002690;
    assign coff[1140] = 256'h00007ae8ffffdc41ffffdc41ffff8518ffff8518000023bf000023bf00007ae8;
    assign coff[1141] = 256'h00003da2ffff8fd1ffff8fd1ffffc25effffc25e0000702f0000702f00003da2;
    assign coff[1142] = 256'h000063dfffffaff1ffffaff1ffff9c21ffff9c210000500f0000500f000063df;
    assign coff[1143] = 256'h00000e03ffff80c5ffff80c5fffff1fdfffff1fd00007f3b00007f3b00000e03;
    assign coff[1144] = 256'h00007dd2ffffe879ffffe879ffff822effff822e000017870000178700007dd2;
    assign coff[1145] = 256'h00004855ffff9666ffff9666ffffb7abffffb7ab0000699a0000699a00004855;
    assign coff[1146] = 256'h00006b3dffffba1effffba1effff94c3ffff94c3000045e2000045e200006b3d;
    assign coff[1147] = 256'h00001a6affff82c1ffff82c1ffffe596ffffe59600007d3f00007d3f00001a6a;
    assign coff[1148] = 256'h000076d0ffffd061ffffd061ffff8930ffff893000002f9f00002f9f000076d0;
    assign coff[1149] = 256'h00003257ffff8a51ffff8a51ffffcda9ffffcda9000075af000075af00003257;
    assign coff[1150] = 256'h00005b8cffffa68affffa68affffa474ffffa474000059760000597600005b8c;
    assign coff[1151] = 256'h00000179ffff8002ffff8002fffffe87fffffe8700007ffe00007ffe00000179;
    assign coff[1152] = 256'h00007fffffffff1effffff1effff8001ffff8001000000e2000000e200007fff;
    assign coff[1153] = 256'h000059e2ffffa4deffffa4deffffa61effffa61e00005b2200005b22000059e2;
    assign coff[1154] = 256'h000075eaffffce34ffffce34ffff8a16ffff8a16000031cc000031cc000075ea;
    assign coff[1155] = 256'h0000302affff8968ffff8968ffffcfd6ffffcfd600007698000076980000302a;
    assign coff[1156] = 256'h00007d5dffffe62affffe62affff82a3ffff82a3000019d6000019d600007d5d;
    assign coff[1157] = 256'h00004660ffff9515ffff9515ffffb9a0ffffb9a000006aeb00006aeb00004660;
    assign coff[1158] = 256'h000069efffffb827ffffb827ffff9611ffff9611000047d9000047d9000069ef;
    assign coff[1159] = 256'h0000181bffff824affff824affffe7e5ffffe7e500007db600007db60000181b;
    assign coff[1160] = 256'h00007f4bfffff293fffff293ffff80b5ffff80b500000d6d00000d6d00007f4b;
    assign coff[1161] = 256'h00005084ffff9c7fffff9c7fffffaf7cffffaf7c000063810000638100005084;
    assign coff[1162] = 256'h00007077ffffc2e2ffffc2e2ffff8f89ffff8f8900003d1e00003d1e00007077;
    assign coff[1163] = 256'h0000244fffff8542ffff8542ffffdbb1ffffdbb100007abe00007abe0000244f;
    assign coff[1164] = 256'h00007a3bffffda00ffffda00ffff85c5ffff85c5000026000000260000007a3b;
    assign coff[1165] = 256'h00003b8fffff8eb3ffff8eb3ffffc471ffffc4710000714d0000714d00003b8f;
    assign coff[1166] = 256'h00006262ffffae1effffae1effff9d9effff9d9e000051e2000051e200006262;
    assign coff[1167] = 256'h00000babffff8088ffff8088fffff455fffff45500007f7800007f7800000bab;
    assign coff[1168] = 256'h00007fcdfffff8d6fffff8d6ffff8033ffff80330000072a0000072a00007fcd;
    assign coff[1169] = 256'h0000554effffa091ffffa091ffffaab2ffffaab200005f6f00005f6f0000554e;
    assign coff[1170] = 256'h00007355ffffc87affffc87affff8cabffff8cab000037860000378600007355;
    assign coff[1171] = 256'h00002a4affff8730ffff8730ffffd5b6ffffd5b6000078d0000078d000002a4a;
    assign coff[1172] = 256'h00007bf2ffffe00bffffe00bffff840effff840e00001ff500001ff500007bf2;
    assign coff[1173] = 256'h0000410cffff91c2ffff91c2ffffbef4ffffbef400006e3e00006e3e0000410c;
    assign coff[1174] = 256'h00006648ffffb30bffffb30bffff99b8ffff99b800004cf500004cf500006648;
    assign coff[1175] = 256'h000011e8ffff8142ffff8142ffffee18ffffee1800007ebe00007ebe000011e8;
    assign coff[1176] = 256'h00007e7bffffec58ffffec58ffff8185ffff8185000013a8000013a800007e7b;
    assign coff[1177] = 256'h00004b8affff98aaffff98aaffffb476ffffb476000067560000675600004b8a;
    assign coff[1178] = 256'h00006d55ffffbd70ffffbd70ffff92abffff92ab000042900000429000006d55;
    assign coff[1179] = 256'h00001e3effff83a0ffff83a0ffffe1c2ffffe1c200007c6000007c6000001e3e;
    assign coff[1180] = 256'h00007838ffffd40cffffd40cffff87c8ffff87c800002bf400002bf400007838;
    assign coff[1181] = 256'h000035edffff8beaffff8beaffffca13ffffca130000741600007416000035ed;
    assign coff[1182] = 256'h00005e3fffffa963ffffa963ffffa1c1ffffa1c10000569d0000569d00005e3f;
    assign coff[1183] = 256'h00000566ffff801dffff801dfffffa9afffffa9a00007fe300007fe300000566;
    assign coff[1184] = 256'h00007ff0fffffbfafffffbfaffff8010ffff8010000004060000040600007ff0;
    assign coff[1185] = 256'h0000579fffffa2b0ffffa2b0ffffa861ffffa86100005d5000005d500000579f;
    assign coff[1186] = 256'h000074a8ffffcb53ffffcb53ffff8b58ffff8b58000034ad000034ad000074a8;
    assign coff[1187] = 256'h00002d3effff8843ffff8843ffffd2c2ffffd2c2000077bd000077bd00002d3e;
    assign coff[1188] = 256'h00007cb1ffffe318ffffe318ffff834fffff834f00001ce800001ce800007cb1;
    assign coff[1189] = 256'h000043bbffff9363ffff9363ffffbc45ffffbc4500006c9d00006c9d000043bb;
    assign coff[1190] = 256'h00006824ffffb593ffffb593ffff97dcffff97dc00004a6d00004a6d00006824;
    assign coff[1191] = 256'h00001503ffff81bdffff81bdffffeafdffffeafd00007e4300007e4300001503;
    assign coff[1192] = 256'h00007eedffffef74ffffef74ffff8113ffff81130000108c0000108c00007eed;
    assign coff[1193] = 256'h00004e0dffff9a8dffff9a8dffffb1f3ffffb1f3000065730000657300004e0d;
    assign coff[1194] = 256'h00006eefffffc024ffffc024ffff9111ffff911100003fdc00003fdc00006eef;
    assign coff[1195] = 256'h00002149ffff8467ffff8467ffffdeb7ffffdeb700007b9900007b9900002149;
    assign coff[1196] = 256'h00007942ffffd703ffffd703ffff86beffff86be000028fd000028fd00007942;
    assign coff[1197] = 256'h000038c2ffff8d46ffff8d46ffffc73effffc73e000072ba000072ba000038c2;
    assign coff[1198] = 256'h00006058ffffabbaffffabbaffff9fa8ffff9fa8000054460000544600006058;
    assign coff[1199] = 256'h00000889ffff8049ffff8049fffff777fffff77700007fb700007fb700000889;
    assign coff[1200] = 256'h00007f96fffff5b4fffff5b4ffff806affff806a00000a4c00000a4c00007f96;
    assign coff[1201] = 256'h000052efffff9e81ffff9e81ffffad11ffffad110000617f0000617f000052ef;
    assign coff[1202] = 256'h000071efffffc5a9ffffc5a9ffff8e11ffff8e1100003a5700003a57000071ef;
    assign coff[1203] = 256'h00002750ffff8630ffff8630ffffd8b0ffffd8b0000079d0000079d000002750;
    assign coff[1204] = 256'h00007b20ffffdd03ffffdd03ffff84e0ffff84e0000022fd000022fd00007b20;
    assign coff[1205] = 256'h00003e52ffff9032ffff9032ffffc1aeffffc1ae00006fce00006fce00003e52;
    assign coff[1206] = 256'h0000645dffffb08effffb08effff9ba3ffff9ba300004f7200004f720000645d;
    assign coff[1207] = 256'h00000ecbffff80dcffff80dcfffff135fffff13500007f2400007f2400000ecb;
    assign coff[1208] = 256'h00007df6ffffe93fffffe93fffff820affff820a000016c1000016c100007df6;
    assign coff[1209] = 256'h000048fbffff96d8ffff96d8ffffb705ffffb7050000692800006928000048fb;
    assign coff[1210] = 256'h00006baaffffbac7ffffbac7ffff9456ffff9456000045390000453900006baa;
    assign coff[1211] = 256'h00001b2fffff82ebffff82ebffffe4d1ffffe4d100007d1500007d1500001b2f;
    assign coff[1212] = 256'h0000771affffd11cffffd11cffff88e6ffff88e600002ee400002ee40000771a;
    assign coff[1213] = 256'h00003310ffff8aa0ffff8aa0ffffccf0ffffccf0000075600000756000003310;
    assign coff[1214] = 256'h00005c18ffffa71affffa71affffa3e8ffffa3e8000058e6000058e600005c18;
    assign coff[1215] = 256'h00000242ffff8005ffff8005fffffdbefffffdbe00007ffb00007ffb00000242;
    assign coff[1216] = 256'h00007ffafffffd8cfffffd8cffff8006ffff8006000002740000027400007ffa;
    assign coff[1217] = 256'h000058c2ffffa3c6ffffa3c6ffffa73effffa73e00005c3a00005c3a000058c2;
    assign coff[1218] = 256'h0000754cffffccc2ffffccc2ffff8ab4ffff8ab40000333e0000333e0000754c;
    assign coff[1219] = 256'h00002eb5ffff88d3ffff88d3ffffd14bffffd14b0000772d0000772d00002eb5;
    assign coff[1220] = 256'h00007d0affffe4a0ffffe4a0ffff82f6ffff82f600001b6000001b6000007d0a;
    assign coff[1221] = 256'h0000450fffff943affff943affffbaf1ffffbaf100006bc600006bc60000450f;
    assign coff[1222] = 256'h0000690cffffb6dcffffb6dcffff96f4ffff96f400004924000049240000690c;
    assign coff[1223] = 256'h0000168fffff8201ffff8201ffffe971ffffe97100007dff00007dff0000168f;
    assign coff[1224] = 256'h00007f1ffffff104fffff104ffff80e1ffff80e100000efc00000efc00007f1f;
    assign coff[1225] = 256'h00004f4affff9b84ffff9b84ffffb0b6ffffb0b60000647c0000647c00004f4a;
    assign coff[1226] = 256'h00006fb5ffffc182ffffc182ffff904bffff904b00003e7e00003e7e00006fb5;
    assign coff[1227] = 256'h000022cdffff84d2ffff84d2ffffdd33ffffdd3300007b2e00007b2e000022cd;
    assign coff[1228] = 256'h000079c1ffffd880ffffd880ffff863fffff863f0000278000002780000079c1;
    assign coff[1229] = 256'h00003a2affff8dfaffff8dfaffffc5d6ffffc5d6000072060000720600003a2a;
    assign coff[1230] = 256'h0000615fffffaceaffffaceaffff9ea1ffff9ea100005316000053160000615f;
    assign coff[1231] = 256'h00000a1affff8066ffff8066fffff5e6fffff5e600007f9a00007f9a00000a1a;
    assign coff[1232] = 256'h00007fb4fffff745fffff745ffff804cffff804c000008bb000008bb00007fb4;
    assign coff[1233] = 256'h00005420ffff9f87ffff9f87ffffabe0ffffabe0000060790000607900005420;
    assign coff[1234] = 256'h000072a4ffffc710ffffc710ffff8d5cffff8d5c000038f0000038f0000072a4;
    assign coff[1235] = 256'h000028ceffff86adffff86adffffd732ffffd7320000795300007953000028ce;
    assign coff[1236] = 256'h00007b8bffffde86ffffde86ffff8475ffff84750000217a0000217a00007b8b;
    assign coff[1237] = 256'h00003fb0ffff90f8ffff90f8ffffc050ffffc05000006f0800006f0800003fb0;
    assign coff[1238] = 256'h00006554ffffb1cbffffb1cbffff9aacffff9aac00004e3500004e3500006554;
    assign coff[1239] = 256'h0000105affff810cffff810cffffefa6ffffefa600007ef400007ef40000105a;
    assign coff[1240] = 256'h00007e3bffffeacbffffeacbffff81c5ffff81c5000015350000153500007e3b;
    assign coff[1241] = 256'h00004a44ffff97bfffff97bfffffb5bcffffb5bc000068410000684100004a44;
    assign coff[1242] = 256'h00006c82ffffbc1affffbc1affff937effff937e000043e6000043e600006c82;
    assign coff[1243] = 256'h00001cb7ffff8343ffff8343ffffe349ffffe34900007cbd00007cbd00001cb7;
    assign coff[1244] = 256'h000077abffffd293ffffd293ffff8855ffff885500002d6d00002d6d000077ab;
    assign coff[1245] = 256'h00003480ffff8b43ffff8b43ffffcb80ffffcb80000074bd000074bd00003480;
    assign coff[1246] = 256'h00005d2dffffa83dffffa83dffffa2d3ffffa2d3000057c3000057c300005d2d;
    assign coff[1247] = 256'h000003d4ffff800fffff800ffffffc2cfffffc2c00007ff100007ff1000003d4;
    assign coff[1248] = 256'h00007fe1fffffa68fffffa68ffff801fffff801f000005980000059800007fe1;
    assign coff[1249] = 256'h00005678ffffa19fffffa19fffffa988ffffa98800005e6100005e6100005678;
    assign coff[1250] = 256'h00007401ffffc9e5ffffc9e5ffff8bffffff8bff0000361b0000361b00007401;
    assign coff[1251] = 256'h00002bc5ffff87b7ffff87b7ffffd43bffffd43b000078490000784900002bc5;
    assign coff[1252] = 256'h00007c54ffffe191ffffe191ffff83acffff83ac00001e6f00001e6f00007c54;
    assign coff[1253] = 256'h00004265ffff9291ffff9291ffffbd9bffffbd9b00006d6f00006d6f00004265;
    assign coff[1254] = 256'h00006738ffffb44effffb44effff98c8ffff98c800004bb200004bb200006738;
    assign coff[1255] = 256'h00001376ffff817dffff817dffffec8affffec8a00007e8300007e8300001376;
    assign coff[1256] = 256'h00007eb7ffffede6ffffede6ffff8149ffff81490000121a0000121a00007eb7;
    assign coff[1257] = 256'h00004ccdffff999affff999affffb333ffffb333000066660000666600004ccd;
    assign coff[1258] = 256'h00006e24ffffbec9ffffbec9ffff91dcffff91dc000041370000413700006e24;
    assign coff[1259] = 256'h00001fc5ffff8401ffff8401ffffe03bffffe03b00007bff00007bff00001fc5;
    assign coff[1260] = 256'h000078bfffffd587ffffd587ffff8741ffff874100002a7900002a79000078bf;
    assign coff[1261] = 256'h00003759ffff8c96ffff8c96ffffc8a7ffffc8a70000736a0000736a00003759;
    assign coff[1262] = 256'h00005f4dffffaa8dffffaa8dffffa0b3ffffa0b3000055730000557300005f4d;
    assign coff[1263] = 256'h000006f8ffff8031ffff8031fffff908fffff90800007fcf00007fcf000006f8;
    assign coff[1264] = 256'h00007f73fffff423fffff423ffff808dffff808d00000bdd00000bdd00007f73;
    assign coff[1265] = 256'h000051bbffff9d7effff9d7effffae45ffffae450000628200006282000051bb;
    assign coff[1266] = 256'h00007135ffffc445ffffc445ffff8ecbffff8ecb00003bbb00003bbb00007135;
    assign coff[1267] = 256'h000025d0ffff85b7ffff85b7ffffda30ffffda3000007a4900007a49000025d0;
    assign coff[1268] = 256'h00007ab0ffffdb80ffffdb80ffff8550ffff8550000024800000248000007ab0;
    assign coff[1269] = 256'h00003cf2ffff8f71ffff8f71ffffc30effffc30e0000708f0000708f00003cf2;
    assign coff[1270] = 256'h00006361ffffaf54ffffaf54ffff9c9fffff9c9f000050ac000050ac00006361;
    assign coff[1271] = 256'h00000d3bffff80b0ffff80b0fffff2c5fffff2c500007f5000007f5000000d3b;
    assign coff[1272] = 256'h00007dacffffe7b4ffffe7b4ffff8254ffff82540000184c0000184c00007dac;
    assign coff[1273] = 256'h000047afffff95f5ffff95f5ffffb851ffffb85100006a0b00006a0b000047af;
    assign coff[1274] = 256'h00006acfffffb976ffffb976ffff9531ffff95310000468a0000468a00006acf;
    assign coff[1275] = 256'h000019a5ffff8298ffff8298ffffe65bffffe65b00007d6800007d68000019a5;
    assign coff[1276] = 256'h00007685ffffcfa7ffffcfa7ffff897bffff897b000030590000305900007685;
    assign coff[1277] = 256'h0000319effff8a02ffff8a02ffffce62ffffce62000075fe000075fe0000319e;
    assign coff[1278] = 256'h00005affffffa5faffffa5faffffa501ffffa50100005a0600005a0600005aff;
    assign coff[1279] = 256'h000000b0ffff8001ffff8001ffffff50ffffff5000007fff00007fff000000b0;
    assign coff[1280] = 256'h00007fffffffff82ffffff82ffff8001ffff80010000007e0000007e00007fff;
    assign coff[1281] = 256'h00005a29ffffa525ffffa525ffffa5d7ffffa5d700005adb00005adb00005a29;
    assign coff[1282] = 256'h00007611ffffce90ffffce90ffff89efffff89ef000031700000317000007611;
    assign coff[1283] = 256'h00003088ffff898effff898effffcf78ffffcf78000076720000767200003088;
    assign coff[1284] = 256'h00007d72ffffe68cffffe68cffff828effff828e000019740000197400007d72;
    assign coff[1285] = 256'h000046b4ffff954dffff954dffffb94cffffb94c00006ab300006ab3000046b4;
    assign coff[1286] = 256'h00006a28ffffb87bffffb87bffff95d8ffff95d8000047850000478500006a28;
    assign coff[1287] = 256'h0000187dffff825dffff825dffffe783ffffe78300007da300007da30000187d;
    assign coff[1288] = 256'h00007f56fffff2f7fffff2f7ffff80aaffff80aa00000d0900000d0900007f56;
    assign coff[1289] = 256'h000050d3ffff9cbeffff9cbeffffaf2dffffaf2d0000634200006342000050d3;
    assign coff[1290] = 256'h000070a7ffffc33bffffc33bffff8f59ffff8f5900003cc500003cc5000070a7;
    assign coff[1291] = 256'h000024b0ffff855fffff855fffffdb50ffffdb5000007aa100007aa1000024b0;
    assign coff[1292] = 256'h00007a58ffffda60ffffda60ffff85a8ffff85a8000025a0000025a000007a58;
    assign coff[1293] = 256'h00003be8ffff8ee2ffff8ee2ffffc418ffffc4180000711e0000711e00003be8;
    assign coff[1294] = 256'h000062a2ffffae6bffffae6bffff9d5effff9d5e0000519500005195000062a2;
    assign coff[1295] = 256'h00000c0fffff8092ffff8092fffff3f1fffff3f100007f6e00007f6e00000c0f;
    assign coff[1296] = 256'h00007fd2fffff93bfffff93bffff802effff802e000006c5000006c500007fd2;
    assign coff[1297] = 256'h00005598ffffa0d4ffffa0d4ffffaa68ffffaa6800005f2c00005f2c00005598;
    assign coff[1298] = 256'h00007380ffffc8d4ffffc8d4ffff8c80ffff8c800000372c0000372c00007380;
    assign coff[1299] = 256'h00002aa9ffff8751ffff8751ffffd557ffffd557000078af000078af00002aa9;
    assign coff[1300] = 256'h00007c0bffffe06cffffe06cffff83f5ffff83f500001f9400001f9400007c0b;
    assign coff[1301] = 256'h00004162ffff91f6ffff91f6ffffbe9effffbe9e00006e0a00006e0a00004162;
    assign coff[1302] = 256'h00006684ffffb35bffffb35bffff997cffff997c00004ca500004ca500006684;
    assign coff[1303] = 256'h0000124cffff8150ffff8150ffffedb4ffffedb400007eb000007eb00000124c;
    assign coff[1304] = 256'h00007e8bffffecbcffffecbcffff8175ffff8175000013440000134400007e8b;
    assign coff[1305] = 256'h00004bdbffff98e6ffff98e6ffffb425ffffb4250000671a0000671a00004bdb;
    assign coff[1306] = 256'h00006d89ffffbdc6ffffbdc6ffff9277ffff92770000423a0000423a00006d89;
    assign coff[1307] = 256'h00001ea0ffff83b8ffff83b8ffffe160ffffe16000007c4800007c4800001ea0;
    assign coff[1308] = 256'h0000785affffd46bffffd46bffff87a6ffff87a600002b9500002b950000785a;
    assign coff[1309] = 256'h00003648ffff8c15ffff8c15ffffc9b8ffffc9b8000073eb000073eb00003648;
    assign coff[1310] = 256'h00005e83ffffa9adffffa9adffffa17dffffa17d000056530000565300005e83;
    assign coff[1311] = 256'h000005caffff8022ffff8022fffffa36fffffa3600007fde00007fde000005ca;
    assign coff[1312] = 256'h00007ff3fffffc5efffffc5effff800dffff800d000003a2000003a200007ff3;
    assign coff[1313] = 256'h000057e8ffffa2f5ffffa2f5ffffa818ffffa81800005d0b00005d0b000057e8;
    assign coff[1314] = 256'h000074d2ffffcbaeffffcbaeffff8b2effff8b2e0000345200003452000074d2;
    assign coff[1315] = 256'h00002d9cffff8867ffff8867ffffd264ffffd264000077990000779900002d9c;
    assign coff[1316] = 256'h00007cc8ffffe37affffe37affff8338ffff833800001c8600001c8600007cc8;
    assign coff[1317] = 256'h00004411ffff9399ffff9399ffffbbefffffbbef00006c6700006c6700004411;
    assign coff[1318] = 256'h0000685effffb5e5ffffb5e5ffff97a2ffff97a200004a1b00004a1b0000685e;
    assign coff[1319] = 256'h00001566ffff81cdffff81cdffffea9affffea9a00007e3300007e3300001566;
    assign coff[1320] = 256'h00007efaffffefd8ffffefd8ffff8106ffff8106000010280000102800007efa;
    assign coff[1321] = 256'h00004e5dffff9acaffff9acaffffb1a3ffffb1a3000065360000653600004e5d;
    assign coff[1322] = 256'h00006f21ffffc07bffffc07bffff90dfffff90df00003f8500003f8500006f21;
    assign coff[1323] = 256'h000021aaffff8482ffff8482ffffde56ffffde5600007b7e00007b7e000021aa;
    assign coff[1324] = 256'h00007962ffffd762ffffd762ffff869effff869e0000289e0000289e00007962;
    assign coff[1325] = 256'h0000391dffff8d73ffff8d73ffffc6e3ffffc6e30000728d0000728d0000391d;
    assign coff[1326] = 256'h0000609affffac06ffffac06ffff9f66ffff9f66000053fa000053fa0000609a;
    assign coff[1327] = 256'h000008edffff8050ffff8050fffff713fffff71300007fb000007fb0000008ed;
    assign coff[1328] = 256'h00007f9efffff618fffff618ffff8062ffff8062000009e8000009e800007f9e;
    assign coff[1329] = 256'h0000533cffff9ec2ffff9ec2ffffacc4ffffacc40000613e0000613e0000533c;
    assign coff[1330] = 256'h0000721cffffc603ffffc603ffff8de4ffff8de4000039fd000039fd0000721c;
    assign coff[1331] = 256'h000027afffff864fffff864fffffd851ffffd851000079b1000079b1000027af;
    assign coff[1332] = 256'h00007b3bffffdd63ffffdd63ffff84c5ffff84c50000229d0000229d00007b3b;
    assign coff[1333] = 256'h00003eaaffff9063ffff9063ffffc156ffffc15600006f9d00006f9d00003eaa;
    assign coff[1334] = 256'h0000649bffffb0ddffffb0ddffff9b65ffff9b6500004f2300004f230000649b;
    assign coff[1335] = 256'h00000f2effff80e7ffff80e7fffff0d2fffff0d200007f1900007f1900000f2e;
    assign coff[1336] = 256'h00007e08ffffe9a2ffffe9a2ffff81f8ffff81f80000165e0000165e00007e08;
    assign coff[1337] = 256'h0000494dffff9711ffff9711ffffb6b3ffffb6b3000068ef000068ef0000494d;
    assign coff[1338] = 256'h00006be1ffffbb1bffffbb1bffff941fffff941f000044e5000044e500006be1;
    assign coff[1339] = 256'h00001b91ffff8301ffff8301ffffe46fffffe46f00007cff00007cff00001b91;
    assign coff[1340] = 256'h0000773fffffd17affffd17affff88c1ffff88c100002e8600002e860000773f;
    assign coff[1341] = 256'h0000336cffff8ac8ffff8ac8ffffcc94ffffcc9400007538000075380000336c;
    assign coff[1342] = 256'h00005c5dffffa762ffffa762ffffa3a3ffffa3a30000589e0000589e00005c5d;
    assign coff[1343] = 256'h000002a7ffff8007ffff8007fffffd59fffffd5900007ff900007ff9000002a7;
    assign coff[1344] = 256'h00007ffcfffffdf0fffffdf0ffff8004ffff8004000002100000021000007ffc;
    assign coff[1345] = 256'h0000590affffa40bffffa40bffffa6f6ffffa6f600005bf500005bf50000590a;
    assign coff[1346] = 256'h00007574ffffcd1effffcd1effff8a8cffff8a8c000032e2000032e200007574;
    assign coff[1347] = 256'h00002f13ffff88f8ffff88f8ffffd0edffffd0ed000077080000770800002f13;
    assign coff[1348] = 256'h00007d1fffffe502ffffe502ffff82e1ffff82e100001afe00001afe00007d1f;
    assign coff[1349] = 256'h00004564ffff9471ffff9471ffffba9cffffba9c00006b8f00006b8f00004564;
    assign coff[1350] = 256'h00006945ffffb72fffffb72fffff96bbffff96bb000048d1000048d100006945;
    assign coff[1351] = 256'h000016f2ffff8213ffff8213ffffe90effffe90e00007ded00007ded000016f2;
    assign coff[1352] = 256'h00007f2afffff167fffff167ffff80d6ffff80d600000e9900000e9900007f2a;
    assign coff[1353] = 256'h00004f99ffff9bc2ffff9bc2ffffb067ffffb0670000643e0000643e00004f99;
    assign coff[1354] = 256'h00006fe6ffffc1daffffc1daffff901affff901a00003e2600003e2600006fe6;
    assign coff[1355] = 256'h0000232effff84eeffff84eeffffdcd2ffffdcd200007b1200007b120000232e;
    assign coff[1356] = 256'h000079e0ffffd8e0ffffd8e0ffff8620ffff86200000272000002720000079e0;
    assign coff[1357] = 256'h00003a83ffff8e28ffff8e28ffffc57dffffc57d000071d8000071d800003a83;
    assign coff[1358] = 256'h000061a0ffffad37ffffad37ffff9e60ffff9e60000052c9000052c9000061a0;
    assign coff[1359] = 256'h00000a7effff806effff806efffff582fffff58200007f9200007f9200000a7e;
    assign coff[1360] = 256'h00007fbafffff7a9fffff7a9ffff8046ffff8046000008570000085700007fba;
    assign coff[1361] = 256'h0000546cffff9fc9ffff9fc9ffffab94ffffab9400006037000060370000546c;
    assign coff[1362] = 256'h000072d0ffffc76bffffc76bffff8d30ffff8d300000389500003895000072d0;
    assign coff[1363] = 256'h0000292dffff86ceffff86ceffffd6d3ffffd6d300007932000079320000292d;
    assign coff[1364] = 256'h00007ba6ffffdee7ffffdee7ffff845affff845a000021190000211900007ba6;
    assign coff[1365] = 256'h00004007ffff912affff912affffbff9ffffbff900006ed600006ed600004007;
    assign coff[1366] = 256'h00006592ffffb21bffffb21bffff9a6effff9a6e00004de500004de500006592;
    assign coff[1367] = 256'h000010bdffff8119ffff8119ffffef43ffffef4300007ee700007ee7000010bd;
    assign coff[1368] = 256'h00007e4cffffeb2fffffeb2fffff81b4ffff81b4000014d1000014d100007e4c;
    assign coff[1369] = 256'h00004a95ffff97faffff97faffffb56bffffb56b000068060000680600004a95;
    assign coff[1370] = 256'h00006cb7ffffbc6fffffbc6fffff9349ffff9349000043910000439100006cb7;
    assign coff[1371] = 256'h00001d19ffff835affff835affffe2e7ffffe2e700007ca600007ca600001d19;
    assign coff[1372] = 256'h000077cfffffd2f1ffffd2f1ffff8831ffff883100002d0f00002d0f000077cf;
    assign coff[1373] = 256'h000034dbffff8b6cffff8b6cffffcb25ffffcb250000749400007494000034db;
    assign coff[1374] = 256'h00005d72ffffa886ffffa886ffffa28effffa28e0000577a0000577a00005d72;
    assign coff[1375] = 256'h00000439ffff8012ffff8012fffffbc7fffffbc700007fee00007fee00000439;
    assign coff[1376] = 256'h00007fe5fffffaccfffffaccffff801bffff801b000005340000053400007fe5;
    assign coff[1377] = 256'h000056c2ffffa1e3ffffa1e3ffffa93effffa93e00005e1d00005e1d000056c2;
    assign coff[1378] = 256'h0000742bffffca40ffffca40ffff8bd5ffff8bd5000035c0000035c00000742b;
    assign coff[1379] = 256'h00002c23ffff87daffff87daffffd3ddffffd3dd000078260000782600002c23;
    assign coff[1380] = 256'h00007c6cffffe1f2ffffe1f2ffff8394ffff839400001e0e00001e0e00007c6c;
    assign coff[1381] = 256'h000042bbffff92c5ffff92c5ffffbd45ffffbd4500006d3b00006d3b000042bb;
    assign coff[1382] = 256'h00006773ffffb49fffffb49fffff988dffff988d00004b6100004b6100006773;
    assign coff[1383] = 256'h000013d9ffff818cffff818cffffec27ffffec2700007e7400007e74000013d9;
    assign coff[1384] = 256'h00007ec5ffffee4affffee4affff813bffff813b000011b6000011b600007ec5;
    assign coff[1385] = 256'h00004d1dffff99d6ffff99d6ffffb2e3ffffb2e30000662a0000662a00004d1d;
    assign coff[1386] = 256'h00006e57ffffbf20ffffbf20ffff91a9ffff91a9000040e0000040e000006e57;
    assign coff[1387] = 256'h00002026ffff841affff841affffdfdaffffdfda00007be600007be600002026;
    assign coff[1388] = 256'h000078e1ffffd5e5ffffd5e5ffff871fffff871f00002a1b00002a1b000078e1;
    assign coff[1389] = 256'h000037b4ffff8cc1ffff8cc1ffffc84cffffc84c0000733f0000733f000037b4;
    assign coff[1390] = 256'h00005f90ffffaad8ffffaad8ffffa070ffffa070000055280000552800005f90;
    assign coff[1391] = 256'h0000075cffff8036ffff8036fffff8a4fffff8a400007fca00007fca0000075c;
    assign coff[1392] = 256'h00007f7cfffff487fffff487ffff8084ffff808400000b7900000b7900007f7c;
    assign coff[1393] = 256'h00005209ffff9dbeffff9dbeffffadf7ffffadf7000062420000624200005209;
    assign coff[1394] = 256'h00007164ffffc49effffc49effff8e9cffff8e9c00003b6200003b6200007164;
    assign coff[1395] = 256'h00002630ffff85d4ffff85d4ffffd9d0ffffd9d000007a2c00007a2c00002630;
    assign coff[1396] = 256'h00007accffffdbe1ffffdbe1ffff8534ffff85340000241f0000241f00007acc;
    assign coff[1397] = 256'h00003d4affff8fa1ffff8fa1ffffc2b6ffffc2b60000705f0000705f00003d4a;
    assign coff[1398] = 256'h000063a0ffffafa3ffffafa3ffff9c60ffff9c600000505d0000505d000063a0;
    assign coff[1399] = 256'h00000d9fffff80baffff80bafffff261fffff26100007f4600007f4600000d9f;
    assign coff[1400] = 256'h00007dbfffffe817ffffe817ffff8241ffff8241000017e9000017e900007dbf;
    assign coff[1401] = 256'h00004802ffff962dffff962dffffb7feffffb7fe000069d3000069d300004802;
    assign coff[1402] = 256'h00006b06ffffb9caffffb9caffff94faffff94fa000046360000463600006b06;
    assign coff[1403] = 256'h00001a08ffff82adffff82adffffe5f8ffffe5f800007d5300007d5300001a08;
    assign coff[1404] = 256'h000076aaffffd004ffffd004ffff8956ffff895600002ffc00002ffc000076aa;
    assign coff[1405] = 256'h000031fbffff8a29ffff8a29ffffce05ffffce05000075d7000075d7000031fb;
    assign coff[1406] = 256'h00005b45ffffa642ffffa642ffffa4bbffffa4bb000059be000059be00005b45;
    assign coff[1407] = 256'h00000114ffff8001ffff8001fffffeecfffffeec00007fff00007fff00000114;
    assign coff[1408] = 256'h00007ffefffffeb9fffffeb9ffff8002ffff8002000001470000014700007ffe;
    assign coff[1409] = 256'h0000599affffa498ffffa498ffffa666ffffa66600005b6800005b680000599a;
    assign coff[1410] = 256'h000075c3ffffcdd7ffffcdd7ffff8a3dffff8a3d0000322900003229000075c3;
    assign coff[1411] = 256'h00002fcdffff8943ffff8943ffffd033ffffd033000076bd000076bd00002fcd;
    assign coff[1412] = 256'h00007d49ffffe5c7ffffe5c7ffff82b7ffff82b700001a3900001a3900007d49;
    assign coff[1413] = 256'h0000460cffff94deffff94deffffb9f4ffffb9f400006b2200006b220000460c;
    assign coff[1414] = 256'h000069b7ffffb7d4ffffb7d4ffff9649ffff96490000482c0000482c000069b7;
    assign coff[1415] = 256'h000017b8ffff8237ffff8237ffffe848ffffe84800007dc900007dc9000017b8;
    assign coff[1416] = 256'h00007f41fffff22ffffff22fffff80bfffff80bf00000dd100000dd100007f41;
    assign coff[1417] = 256'h00005036ffff9c40ffff9c40ffffafcaffffafca000063c0000063c000005036;
    assign coff[1418] = 256'h00007047ffffc28affffc28affff8fb9ffff8fb900003d7600003d7600007047;
    assign coff[1419] = 256'h000023efffff8526ffff8526ffffdc11ffffdc1100007ada00007ada000023ef;
    assign coff[1420] = 256'h00007a1dffffd9a0ffffd9a0ffff85e3ffff85e3000026600000266000007a1d;
    assign coff[1421] = 256'h00003b36ffff8e85ffff8e85ffffc4caffffc4ca0000717b0000717b00003b36;
    assign coff[1422] = 256'h00006221ffffadd1ffffadd1ffff9ddfffff9ddf0000522f0000522f00006221;
    assign coff[1423] = 256'h00000b47ffff807fffff807ffffff4b9fffff4b900007f8100007f8100000b47;
    assign coff[1424] = 256'h00007fc7fffff872fffff872ffff8039ffff80390000078e0000078e00007fc7;
    assign coff[1425] = 256'h00005502ffffa04effffa04effffaafeffffaafe00005fb200005fb200005502;
    assign coff[1426] = 256'h00007329ffffc81fffffc81fffff8cd7ffff8cd7000037e1000037e100007329;
    assign coff[1427] = 256'h000029ebffff870fffff870fffffd615ffffd615000078f1000078f1000029eb;
    assign coff[1428] = 256'h00007bd9ffffdfa9ffffdfa9ffff8427ffff8427000020570000205700007bd9;
    assign coff[1429] = 256'h000040b5ffff918fffff918fffffbf4bffffbf4b00006e7100006e71000040b5;
    assign coff[1430] = 256'h0000660cffffb2bbffffb2bbffff99f4ffff99f400004d4500004d450000660c;
    assign coff[1431] = 256'h00001185ffff8134ffff8134ffffee7bffffee7b00007ecc00007ecc00001185;
    assign coff[1432] = 256'h00007e6cffffebf5ffffebf5ffff8194ffff81940000140b0000140b00007e6c;
    assign coff[1433] = 256'h00004b38ffff986fffff986fffffb4c8ffffb4c8000067910000679100004b38;
    assign coff[1434] = 256'h00006d21ffffbd1affffbd1affff92dfffff92df000042e6000042e600006d21;
    assign coff[1435] = 256'h00001dddffff8388ffff8388ffffe223ffffe22300007c7800007c7800001ddd;
    assign coff[1436] = 256'h00007815ffffd3aeffffd3aeffff87ebffff87eb00002c5200002c5200007815;
    assign coff[1437] = 256'h00003592ffff8bc0ffff8bc0ffffca6effffca6e000074400000744000003592;
    assign coff[1438] = 256'h00005dfbffffa919ffffa919ffffa205ffffa205000056e7000056e700005dfb;
    assign coff[1439] = 256'h00000501ffff8019ffff8019fffffafffffffaff00007fe700007fe700000501;
    assign coff[1440] = 256'h00007fecfffffb95fffffb95ffff8014ffff80140000046b0000046b00007fec;
    assign coff[1441] = 256'h00005755ffffa26cffffa26cffffa8abffffa8ab00005d9400005d9400005755;
    assign coff[1442] = 256'h0000747fffffcaf7ffffcaf7ffff8b81ffff8b8100003509000035090000747f;
    assign coff[1443] = 256'h00002ce0ffff8820ffff8820ffffd320ffffd320000077e0000077e000002ce0;
    assign coff[1444] = 256'h00007c9bffffe2b6ffffe2b6ffff8365ffff836500001d4a00001d4a00007c9b;
    assign coff[1445] = 256'h00004366ffff932effff932effffbc9affffbc9a00006cd200006cd200004366;
    assign coff[1446] = 256'h000067e9ffffb542ffffb542ffff9817ffff981700004abe00004abe000067e9;
    assign coff[1447] = 256'h000014a0ffff81acffff81acffffeb60ffffeb6000007e5400007e54000014a0;
    assign coff[1448] = 256'h00007ee0ffffef11ffffef11ffff8120ffff8120000010ef000010ef00007ee0;
    assign coff[1449] = 256'h00004dbdffff9a50ffff9a50ffffb243ffffb243000065b0000065b000004dbd;
    assign coff[1450] = 256'h00006ebdffffbfcdffffbfcdffff9143ffff9143000040330000403300006ebd;
    assign coff[1451] = 256'h000020e8ffff844dffff844dffffdf18ffffdf1800007bb300007bb3000020e8;
    assign coff[1452] = 256'h00007922ffffd6a4ffffd6a4ffff86deffff86de0000295c0000295c00007922;
    assign coff[1453] = 256'h00003868ffff8d19ffff8d19ffffc798ffffc798000072e7000072e700003868;
    assign coff[1454] = 256'h00006016ffffab6fffffab6fffff9feaffff9fea000054910000549100006016;
    assign coff[1455] = 256'h00000825ffff8042ffff8042fffff7dbfffff7db00007fbe00007fbe00000825;
    assign coff[1456] = 256'h00007f8efffff550fffff550ffff8072ffff807200000ab000000ab000007f8e;
    assign coff[1457] = 256'h000052a3ffff9e40ffff9e40ffffad5dffffad5d000061c0000061c0000052a3;
    assign coff[1458] = 256'h000071c1ffffc550ffffc550ffff8e3fffff8e3f00003ab000003ab0000071c1;
    assign coff[1459] = 256'h000026f0ffff8611ffff8611ffffd910ffffd910000079ef000079ef000026f0;
    assign coff[1460] = 256'h00007b04ffffdca2ffffdca2ffff84fcffff84fc0000235e0000235e00007b04;
    assign coff[1461] = 256'h00003dfaffff9001ffff9001ffffc206ffffc20600006fff00006fff00003dfa;
    assign coff[1462] = 256'h0000641effffb040ffffb040ffff9be2ffff9be200004fc000004fc00000641e;
    assign coff[1463] = 256'h00000e67ffff80d0ffff80d0fffff199fffff19900007f3000007f3000000e67;
    assign coff[1464] = 256'h00007de4ffffe8dcffffe8dcffff821cffff821c000017240000172400007de4;
    assign coff[1465] = 256'h000048a8ffff969fffff969fffffb758ffffb7580000696100006961000048a8;
    assign coff[1466] = 256'h00006b74ffffba72ffffba72ffff948cffff948c0000458e0000458e00006b74;
    assign coff[1467] = 256'h00001accffff82d6ffff82d6ffffe534ffffe53400007d2a00007d2a00001acc;
    assign coff[1468] = 256'h000076f5ffffd0bfffffd0bfffff890bffff890b00002f4100002f41000076f5;
    assign coff[1469] = 256'h000032b4ffff8a78ffff8a78ffffcd4cffffcd4c0000758800007588000032b4;
    assign coff[1470] = 256'h00005bd2ffffa6d2ffffa6d2ffffa42effffa42e0000592e0000592e00005bd2;
    assign coff[1471] = 256'h000001deffff8003ffff8003fffffe22fffffe2200007ffd00007ffd000001de;
    assign coff[1472] = 256'h00007ff8fffffd27fffffd27ffff8008ffff8008000002d9000002d900007ff8;
    assign coff[1473] = 256'h00005879ffffa380ffffa380ffffa787ffffa78700005c8000005c8000005879;
    assign coff[1474] = 256'h00007523ffffcc66ffffcc66ffff8addffff8add0000339a0000339a00007523;
    assign coff[1475] = 256'h00002e57ffff88afffff88afffffd1a9ffffd1a9000077510000775100002e57;
    assign coff[1476] = 256'h00007cf4ffffe43effffe43effff830cffff830c00001bc200001bc200007cf4;
    assign coff[1477] = 256'h000044baffff9404ffff9404ffffbb46ffffbb4600006bfc00006bfc000044ba;
    assign coff[1478] = 256'h000068d2ffffb68affffb68affff972effff972e0000497600004976000068d2;
    assign coff[1479] = 256'h0000162cffff81efffff81efffffe9d4ffffe9d400007e1100007e110000162c;
    assign coff[1480] = 256'h00007f13fffff0a0fffff0a0ffff80edffff80ed00000f6000000f6000007f13;
    assign coff[1481] = 256'h00004efbffff9b46ffff9b46ffffb105ffffb105000064ba000064ba00004efb;
    assign coff[1482] = 256'h00006f84ffffc12affffc12affff907cffff907c00003ed600003ed600006f84;
    assign coff[1483] = 256'h0000226cffff84b7ffff84b7ffffdd94ffffdd9400007b4900007b490000226c;
    assign coff[1484] = 256'h000079a2ffffd821ffffd821ffff865effff865e000027df000027df000079a2;
    assign coff[1485] = 256'h000039d0ffff8dcdffff8dcdffffc630ffffc6300000723300007233000039d0;
    assign coff[1486] = 256'h0000611dffffac9effffac9effff9ee3ffff9ee300005362000053620000611d;
    assign coff[1487] = 256'h000009b6ffff805effff805efffff64afffff64a00007fa200007fa2000009b6;
    assign coff[1488] = 256'h00007fadfffff6e1fffff6e1ffff8053ffff80530000091f0000091f00007fad;
    assign coff[1489] = 256'h000053d4ffff9f45ffff9f45ffffac2cffffac2c000060bb000060bb000053d4;
    assign coff[1490] = 256'h00007277ffffc6b7ffffc6b7ffff8d89ffff8d89000039490000394900007277;
    assign coff[1491] = 256'h0000286effff868effff868effffd792ffffd79200007972000079720000286e;
    assign coff[1492] = 256'h00007b71ffffde25ffffde25ffff848fffff848f000021db000021db00007b71;
    assign coff[1493] = 256'h00003f59ffff90c6ffff90c6ffffc0a7ffffc0a700006f3a00006f3a00003f59;
    assign coff[1494] = 256'h00006517ffffb17cffffb17cffff9ae9ffff9ae900004e8400004e8400006517;
    assign coff[1495] = 256'h00000ff6ffff8100ffff8100fffff00afffff00a00007f0000007f0000000ff6;
    assign coff[1496] = 256'h00007e2affffea68ffffea68ffff81d6ffff81d6000015980000159800007e2a;
    assign coff[1497] = 256'h000049f2ffff9785ffff9785ffffb60effffb60e0000687b0000687b000049f2;
    assign coff[1498] = 256'h00006c4cffffbbc5ffffbbc5ffff93b4ffff93b40000443b0000443b00006c4c;
    assign coff[1499] = 256'h00001c55ffff832dffff832dffffe3abffffe3ab00007cd300007cd300001c55;
    assign coff[1500] = 256'h00007787ffffd235ffffd235ffff8879ffff887900002dcb00002dcb00007787;
    assign coff[1501] = 256'h00003424ffff8b1affff8b1affffcbdcffffcbdc000074e6000074e600003424;
    assign coff[1502] = 256'h00005ce8ffffa7f4ffffa7f4ffffa318ffffa3180000580c0000580c00005ce8;
    assign coff[1503] = 256'h00000370ffff800cffff800cfffffc90fffffc9000007ff400007ff400000370;
    assign coff[1504] = 256'h00007fdcfffffa03fffffa03ffff8024ffff8024000005fd000005fd00007fdc;
    assign coff[1505] = 256'h0000562dffffa15bffffa15bffffa9d3ffffa9d300005ea500005ea50000562d;
    assign coff[1506] = 256'h000073d6ffffc98affffc98affff8c2affff8c2a0000367600003676000073d6;
    assign coff[1507] = 256'h00002b66ffff8795ffff8795ffffd49affffd49a0000786b0000786b00002b66;
    assign coff[1508] = 256'h00007c3cffffe12fffffe12fffff83c4ffff83c400001ed100001ed100007c3c;
    assign coff[1509] = 256'h0000420fffff925dffff925dffffbdf1ffffbdf100006da300006da30000420f;
    assign coff[1510] = 256'h000066fcffffb3fdffffb3fdffff9904ffff990400004c0300004c03000066fc;
    assign coff[1511] = 256'h00001313ffff816effff816effffecedffffeced00007e9200007e9200001313;
    assign coff[1512] = 256'h00007ea8ffffed83ffffed83ffff8158ffff81580000127d0000127d00007ea8;
    assign coff[1513] = 256'h00004c7cffff995dffff995dffffb384ffffb384000066a3000066a300004c7c;
    assign coff[1514] = 256'h00006df1ffffbe73ffffbe73ffff920fffff920f0000418d0000418d00006df1;
    assign coff[1515] = 256'h00001f63ffff83e8ffff83e8ffffe09dffffe09d00007c1800007c1800001f63;
    assign coff[1516] = 256'h0000789effffd528ffffd528ffff8762ffff876200002ad800002ad80000789e;
    assign coff[1517] = 256'h000036feffff8c6affff8c6affffc902ffffc9020000739600007396000036fe;
    assign coff[1518] = 256'h00005f0affffaa42ffffaa42ffffa0f6ffffa0f6000055be000055be00005f0a;
    assign coff[1519] = 256'h00000693ffff802bffff802bfffff96dfffff96d00007fd500007fd500000693;
    assign coff[1520] = 256'h00007f6afffff3bffffff3bfffff8096ffff809600000c4100000c4100007f6a;
    assign coff[1521] = 256'h0000516effff9d3effff9d3effffae92ffffae92000062c2000062c20000516e;
    assign coff[1522] = 256'h00007106ffffc3ecffffc3ecffff8efaffff8efa00003c1400003c1400007106;
    assign coff[1523] = 256'h00002570ffff8599ffff8599ffffda90ffffda9000007a6700007a6700002570;
    assign coff[1524] = 256'h00007a93ffffdb20ffffdb20ffff856dffff856d000024e0000024e000007a93;
    assign coff[1525] = 256'h00003c99ffff8f41ffff8f41ffffc367ffffc367000070bf000070bf00003c99;
    assign coff[1526] = 256'h00006322ffffaf07ffffaf07ffff9cdeffff9cde000050f9000050f900006322;
    assign coff[1527] = 256'h00000cd7ffff80a5ffff80a5fffff329fffff32900007f5b00007f5b00000cd7;
    assign coff[1528] = 256'h00007d99ffffe751ffffe751ffff8267ffff8267000018af000018af00007d99;
    assign coff[1529] = 256'h0000475cffff95bcffff95bcffffb8a4ffffb8a400006a4400006a440000475c;
    assign coff[1530] = 256'h00006a97ffffb922ffffb922ffff9569ffff9569000046de000046de00006a97;
    assign coff[1531] = 256'h00001943ffff8284ffff8284ffffe6bdffffe6bd00007d7c00007d7c00001943;
    assign coff[1532] = 256'h0000765effffcf4affffcf4affff89a2ffff89a2000030b6000030b60000765e;
    assign coff[1533] = 256'h00003141ffff89dbffff89dbffffcebfffffcebf000076250000762500003141;
    assign coff[1534] = 256'h00005ab8ffffa5b3ffffa5b3ffffa548ffffa54800005a4d00005a4d00005ab8;
    assign coff[1535] = 256'h0000004bffff8001ffff8001ffffffb5ffffffb500007fff00007fff0000004b;
    assign coff[1536] = 256'h00007fffffffffb5ffffffb5ffff8001ffff80010000004b0000004b00007fff;
    assign coff[1537] = 256'h00005a4dffffa548ffffa548ffffa5b3ffffa5b300005ab800005ab800005a4d;
    assign coff[1538] = 256'h00007625ffffcebfffffcebfffff89dbffff89db000031410000314100007625;
    assign coff[1539] = 256'h000030b6ffff89a2ffff89a2ffffcf4affffcf4a0000765e0000765e000030b6;
    assign coff[1540] = 256'h00007d7cffffe6bdffffe6bdffff8284ffff8284000019430000194300007d7c;
    assign coff[1541] = 256'h000046deffff9569ffff9569ffffb922ffffb92200006a9700006a97000046de;
    assign coff[1542] = 256'h00006a44ffffb8a4ffffb8a4ffff95bcffff95bc0000475c0000475c00006a44;
    assign coff[1543] = 256'h000018afffff8267ffff8267ffffe751ffffe75100007d9900007d99000018af;
    assign coff[1544] = 256'h00007f5bfffff329fffff329ffff80a5ffff80a500000cd700000cd700007f5b;
    assign coff[1545] = 256'h000050f9ffff9cdeffff9cdeffffaf07ffffaf070000632200006322000050f9;
    assign coff[1546] = 256'h000070bfffffc367ffffc367ffff8f41ffff8f4100003c9900003c99000070bf;
    assign coff[1547] = 256'h000024e0ffff856dffff856dffffdb20ffffdb2000007a9300007a93000024e0;
    assign coff[1548] = 256'h00007a67ffffda90ffffda90ffff8599ffff8599000025700000257000007a67;
    assign coff[1549] = 256'h00003c14ffff8efaffff8efaffffc3ecffffc3ec000071060000710600003c14;
    assign coff[1550] = 256'h000062c2ffffae92ffffae92ffff9d3effff9d3e0000516e0000516e000062c2;
    assign coff[1551] = 256'h00000c41ffff8096ffff8096fffff3bffffff3bf00007f6a00007f6a00000c41;
    assign coff[1552] = 256'h00007fd5fffff96dfffff96dffff802bffff802b000006930000069300007fd5;
    assign coff[1553] = 256'h000055beffffa0f6ffffa0f6ffffaa42ffffaa4200005f0a00005f0a000055be;
    assign coff[1554] = 256'h00007396ffffc902ffffc902ffff8c6affff8c6a000036fe000036fe00007396;
    assign coff[1555] = 256'h00002ad8ffff8762ffff8762ffffd528ffffd5280000789e0000789e00002ad8;
    assign coff[1556] = 256'h00007c18ffffe09dffffe09dffff83e8ffff83e800001f6300001f6300007c18;
    assign coff[1557] = 256'h0000418dffff920fffff920fffffbe73ffffbe7300006df100006df10000418d;
    assign coff[1558] = 256'h000066a3ffffb384ffffb384ffff995dffff995d00004c7c00004c7c000066a3;
    assign coff[1559] = 256'h0000127dffff8158ffff8158ffffed83ffffed8300007ea800007ea80000127d;
    assign coff[1560] = 256'h00007e92ffffecedffffecedffff816effff816e000013130000131300007e92;
    assign coff[1561] = 256'h00004c03ffff9904ffff9904ffffb3fdffffb3fd000066fc000066fc00004c03;
    assign coff[1562] = 256'h00006da3ffffbdf1ffffbdf1ffff925dffff925d0000420f0000420f00006da3;
    assign coff[1563] = 256'h00001ed1ffff83c4ffff83c4ffffe12fffffe12f00007c3c00007c3c00001ed1;
    assign coff[1564] = 256'h0000786bffffd49affffd49affff8795ffff879500002b6600002b660000786b;
    assign coff[1565] = 256'h00003676ffff8c2affff8c2affffc98affffc98a000073d6000073d600003676;
    assign coff[1566] = 256'h00005ea5ffffa9d3ffffa9d3ffffa15bffffa15b0000562d0000562d00005ea5;
    assign coff[1567] = 256'h000005fdffff8024ffff8024fffffa03fffffa0300007fdc00007fdc000005fd;
    assign coff[1568] = 256'h00007ff4fffffc90fffffc90ffff800cffff800c000003700000037000007ff4;
    assign coff[1569] = 256'h0000580cffffa318ffffa318ffffa7f4ffffa7f400005ce800005ce80000580c;
    assign coff[1570] = 256'h000074e6ffffcbdcffffcbdcffff8b1affff8b1a0000342400003424000074e6;
    assign coff[1571] = 256'h00002dcbffff8879ffff8879ffffd235ffffd235000077870000778700002dcb;
    assign coff[1572] = 256'h00007cd3ffffe3abffffe3abffff832dffff832d00001c5500001c5500007cd3;
    assign coff[1573] = 256'h0000443bffff93b4ffff93b4ffffbbc5ffffbbc500006c4c00006c4c0000443b;
    assign coff[1574] = 256'h0000687bffffb60effffb60effff9785ffff9785000049f2000049f20000687b;
    assign coff[1575] = 256'h00001598ffff81d6ffff81d6ffffea68ffffea6800007e2a00007e2a00001598;
    assign coff[1576] = 256'h00007f00fffff00afffff00affff8100ffff810000000ff600000ff600007f00;
    assign coff[1577] = 256'h00004e84ffff9ae9ffff9ae9ffffb17cffffb17c000065170000651700004e84;
    assign coff[1578] = 256'h00006f3affffc0a7ffffc0a7ffff90c6ffff90c600003f5900003f5900006f3a;
    assign coff[1579] = 256'h000021dbffff848fffff848fffffde25ffffde2500007b7100007b71000021db;
    assign coff[1580] = 256'h00007972ffffd792ffffd792ffff868effff868e0000286e0000286e00007972;
    assign coff[1581] = 256'h00003949ffff8d89ffff8d89ffffc6b7ffffc6b7000072770000727700003949;
    assign coff[1582] = 256'h000060bbffffac2cffffac2cffff9f45ffff9f45000053d4000053d4000060bb;
    assign coff[1583] = 256'h0000091fffff8053ffff8053fffff6e1fffff6e100007fad00007fad0000091f;
    assign coff[1584] = 256'h00007fa2fffff64afffff64affff805effff805e000009b6000009b600007fa2;
    assign coff[1585] = 256'h00005362ffff9ee3ffff9ee3ffffac9effffac9e0000611d0000611d00005362;
    assign coff[1586] = 256'h00007233ffffc630ffffc630ffff8dcdffff8dcd000039d0000039d000007233;
    assign coff[1587] = 256'h000027dfffff865effff865effffd821ffffd821000079a2000079a2000027df;
    assign coff[1588] = 256'h00007b49ffffdd94ffffdd94ffff84b7ffff84b70000226c0000226c00007b49;
    assign coff[1589] = 256'h00003ed6ffff907cffff907cffffc12affffc12a00006f8400006f8400003ed6;
    assign coff[1590] = 256'h000064baffffb105ffffb105ffff9b46ffff9b4600004efb00004efb000064ba;
    assign coff[1591] = 256'h00000f60ffff80edffff80edfffff0a0fffff0a000007f1300007f1300000f60;
    assign coff[1592] = 256'h00007e11ffffe9d4ffffe9d4ffff81efffff81ef0000162c0000162c00007e11;
    assign coff[1593] = 256'h00004976ffff972effff972effffb68affffb68a000068d2000068d200004976;
    assign coff[1594] = 256'h00006bfcffffbb46ffffbb46ffff9404ffff9404000044ba000044ba00006bfc;
    assign coff[1595] = 256'h00001bc2ffff830cffff830cffffe43effffe43e00007cf400007cf400001bc2;
    assign coff[1596] = 256'h00007751ffffd1a9ffffd1a9ffff88afffff88af00002e5700002e5700007751;
    assign coff[1597] = 256'h0000339affff8addffff8addffffcc66ffffcc6600007523000075230000339a;
    assign coff[1598] = 256'h00005c80ffffa787ffffa787ffffa380ffffa380000058790000587900005c80;
    assign coff[1599] = 256'h000002d9ffff8008ffff8008fffffd27fffffd2700007ff800007ff8000002d9;
    assign coff[1600] = 256'h00007ffdfffffe22fffffe22ffff8003ffff8003000001de000001de00007ffd;
    assign coff[1601] = 256'h0000592effffa42effffa42effffa6d2ffffa6d200005bd200005bd20000592e;
    assign coff[1602] = 256'h00007588ffffcd4cffffcd4cffff8a78ffff8a78000032b4000032b400007588;
    assign coff[1603] = 256'h00002f41ffff890bffff890bffffd0bfffffd0bf000076f5000076f500002f41;
    assign coff[1604] = 256'h00007d2affffe534ffffe534ffff82d6ffff82d600001acc00001acc00007d2a;
    assign coff[1605] = 256'h0000458effff948cffff948cffffba72ffffba7200006b7400006b740000458e;
    assign coff[1606] = 256'h00006961ffffb758ffffb758ffff969fffff969f000048a8000048a800006961;
    assign coff[1607] = 256'h00001724ffff821cffff821cffffe8dcffffe8dc00007de400007de400001724;
    assign coff[1608] = 256'h00007f30fffff199fffff199ffff80d0ffff80d000000e6700000e6700007f30;
    assign coff[1609] = 256'h00004fc0ffff9be2ffff9be2ffffb040ffffb0400000641e0000641e00004fc0;
    assign coff[1610] = 256'h00006fffffffc206ffffc206ffff9001ffff900100003dfa00003dfa00006fff;
    assign coff[1611] = 256'h0000235effff84fcffff84fcffffdca2ffffdca200007b0400007b040000235e;
    assign coff[1612] = 256'h000079efffffd910ffffd910ffff8611ffff8611000026f0000026f0000079ef;
    assign coff[1613] = 256'h00003ab0ffff8e3fffff8e3fffffc550ffffc550000071c1000071c100003ab0;
    assign coff[1614] = 256'h000061c0ffffad5dffffad5dffff9e40ffff9e40000052a3000052a3000061c0;
    assign coff[1615] = 256'h00000ab0ffff8072ffff8072fffff550fffff55000007f8e00007f8e00000ab0;
    assign coff[1616] = 256'h00007fbefffff7dbfffff7dbffff8042ffff8042000008250000082500007fbe;
    assign coff[1617] = 256'h00005491ffff9feaffff9feaffffab6fffffab6f000060160000601600005491;
    assign coff[1618] = 256'h000072e7ffffc798ffffc798ffff8d19ffff8d190000386800003868000072e7;
    assign coff[1619] = 256'h0000295cffff86deffff86deffffd6a4ffffd6a400007922000079220000295c;
    assign coff[1620] = 256'h00007bb3ffffdf18ffffdf18ffff844dffff844d000020e8000020e800007bb3;
    assign coff[1621] = 256'h00004033ffff9143ffff9143ffffbfcdffffbfcd00006ebd00006ebd00004033;
    assign coff[1622] = 256'h000065b0ffffb243ffffb243ffff9a50ffff9a5000004dbd00004dbd000065b0;
    assign coff[1623] = 256'h000010efffff8120ffff8120ffffef11ffffef1100007ee000007ee0000010ef;
    assign coff[1624] = 256'h00007e54ffffeb60ffffeb60ffff81acffff81ac000014a0000014a000007e54;
    assign coff[1625] = 256'h00004abeffff9817ffff9817ffffb542ffffb542000067e9000067e900004abe;
    assign coff[1626] = 256'h00006cd2ffffbc9affffbc9affff932effff932e000043660000436600006cd2;
    assign coff[1627] = 256'h00001d4affff8365ffff8365ffffe2b6ffffe2b600007c9b00007c9b00001d4a;
    assign coff[1628] = 256'h000077e0ffffd320ffffd320ffff8820ffff882000002ce000002ce0000077e0;
    assign coff[1629] = 256'h00003509ffff8b81ffff8b81ffffcaf7ffffcaf70000747f0000747f00003509;
    assign coff[1630] = 256'h00005d94ffffa8abffffa8abffffa26cffffa26c000057550000575500005d94;
    assign coff[1631] = 256'h0000046bffff8014ffff8014fffffb95fffffb9500007fec00007fec0000046b;
    assign coff[1632] = 256'h00007fe7fffffafffffffaffffff8019ffff8019000005010000050100007fe7;
    assign coff[1633] = 256'h000056e7ffffa205ffffa205ffffa919ffffa91900005dfb00005dfb000056e7;
    assign coff[1634] = 256'h00007440ffffca6effffca6effff8bc0ffff8bc0000035920000359200007440;
    assign coff[1635] = 256'h00002c52ffff87ebffff87ebffffd3aeffffd3ae000078150000781500002c52;
    assign coff[1636] = 256'h00007c78ffffe223ffffe223ffff8388ffff838800001ddd00001ddd00007c78;
    assign coff[1637] = 256'h000042e6ffff92dfffff92dfffffbd1affffbd1a00006d2100006d21000042e6;
    assign coff[1638] = 256'h00006791ffffb4c8ffffb4c8ffff986fffff986f00004b3800004b3800006791;
    assign coff[1639] = 256'h0000140bffff8194ffff8194ffffebf5ffffebf500007e6c00007e6c0000140b;
    assign coff[1640] = 256'h00007eccffffee7bffffee7bffff8134ffff8134000011850000118500007ecc;
    assign coff[1641] = 256'h00004d45ffff99f4ffff99f4ffffb2bbffffb2bb0000660c0000660c00004d45;
    assign coff[1642] = 256'h00006e71ffffbf4bffffbf4bffff918fffff918f000040b5000040b500006e71;
    assign coff[1643] = 256'h00002057ffff8427ffff8427ffffdfa9ffffdfa900007bd900007bd900002057;
    assign coff[1644] = 256'h000078f1ffffd615ffffd615ffff870fffff870f000029eb000029eb000078f1;
    assign coff[1645] = 256'h000037e1ffff8cd7ffff8cd7ffffc81fffffc81f0000732900007329000037e1;
    assign coff[1646] = 256'h00005fb2ffffaafeffffaafeffffa04effffa04e000055020000550200005fb2;
    assign coff[1647] = 256'h0000078effff8039ffff8039fffff872fffff87200007fc700007fc70000078e;
    assign coff[1648] = 256'h00007f81fffff4b9fffff4b9ffff807fffff807f00000b4700000b4700007f81;
    assign coff[1649] = 256'h0000522fffff9ddfffff9ddfffffadd1ffffadd100006221000062210000522f;
    assign coff[1650] = 256'h0000717bffffc4caffffc4caffff8e85ffff8e8500003b3600003b360000717b;
    assign coff[1651] = 256'h00002660ffff85e3ffff85e3ffffd9a0ffffd9a000007a1d00007a1d00002660;
    assign coff[1652] = 256'h00007adaffffdc11ffffdc11ffff8526ffff8526000023ef000023ef00007ada;
    assign coff[1653] = 256'h00003d76ffff8fb9ffff8fb9ffffc28affffc28a000070470000704700003d76;
    assign coff[1654] = 256'h000063c0ffffafcaffffafcaffff9c40ffff9c400000503600005036000063c0;
    assign coff[1655] = 256'h00000dd1ffff80bfffff80bffffff22ffffff22f00007f4100007f4100000dd1;
    assign coff[1656] = 256'h00007dc9ffffe848ffffe848ffff8237ffff8237000017b8000017b800007dc9;
    assign coff[1657] = 256'h0000482cffff9649ffff9649ffffb7d4ffffb7d4000069b7000069b70000482c;
    assign coff[1658] = 256'h00006b22ffffb9f4ffffb9f4ffff94deffff94de0000460c0000460c00006b22;
    assign coff[1659] = 256'h00001a39ffff82b7ffff82b7ffffe5c7ffffe5c700007d4900007d4900001a39;
    assign coff[1660] = 256'h000076bdffffd033ffffd033ffff8943ffff894300002fcd00002fcd000076bd;
    assign coff[1661] = 256'h00003229ffff8a3dffff8a3dffffcdd7ffffcdd7000075c3000075c300003229;
    assign coff[1662] = 256'h00005b68ffffa666ffffa666ffffa498ffffa4980000599a0000599a00005b68;
    assign coff[1663] = 256'h00000147ffff8002ffff8002fffffeb9fffffeb900007ffe00007ffe00000147;
    assign coff[1664] = 256'h00007ffffffffeecfffffeecffff8001ffff8001000001140000011400007fff;
    assign coff[1665] = 256'h000059beffffa4bbffffa4bbffffa642ffffa64200005b4500005b45000059be;
    assign coff[1666] = 256'h000075d7ffffce05ffffce05ffff8a29ffff8a29000031fb000031fb000075d7;
    assign coff[1667] = 256'h00002ffcffff8956ffff8956ffffd004ffffd004000076aa000076aa00002ffc;
    assign coff[1668] = 256'h00007d53ffffe5f8ffffe5f8ffff82adffff82ad00001a0800001a0800007d53;
    assign coff[1669] = 256'h00004636ffff94faffff94faffffb9caffffb9ca00006b0600006b0600004636;
    assign coff[1670] = 256'h000069d3ffffb7feffffb7feffff962dffff962d0000480200004802000069d3;
    assign coff[1671] = 256'h000017e9ffff8241ffff8241ffffe817ffffe81700007dbf00007dbf000017e9;
    assign coff[1672] = 256'h00007f46fffff261fffff261ffff80baffff80ba00000d9f00000d9f00007f46;
    assign coff[1673] = 256'h0000505dffff9c60ffff9c60ffffafa3ffffafa3000063a0000063a00000505d;
    assign coff[1674] = 256'h0000705fffffc2b6ffffc2b6ffff8fa1ffff8fa100003d4a00003d4a0000705f;
    assign coff[1675] = 256'h0000241fffff8534ffff8534ffffdbe1ffffdbe100007acc00007acc0000241f;
    assign coff[1676] = 256'h00007a2cffffd9d0ffffd9d0ffff85d4ffff85d4000026300000263000007a2c;
    assign coff[1677] = 256'h00003b62ffff8e9cffff8e9cffffc49effffc49e000071640000716400003b62;
    assign coff[1678] = 256'h00006242ffffadf7ffffadf7ffff9dbeffff9dbe000052090000520900006242;
    assign coff[1679] = 256'h00000b79ffff8084ffff8084fffff487fffff48700007f7c00007f7c00000b79;
    assign coff[1680] = 256'h00007fcafffff8a4fffff8a4ffff8036ffff80360000075c0000075c00007fca;
    assign coff[1681] = 256'h00005528ffffa070ffffa070ffffaad8ffffaad800005f9000005f9000005528;
    assign coff[1682] = 256'h0000733fffffc84cffffc84cffff8cc1ffff8cc1000037b4000037b40000733f;
    assign coff[1683] = 256'h00002a1bffff871fffff871fffffd5e5ffffd5e5000078e1000078e100002a1b;
    assign coff[1684] = 256'h00007be6ffffdfdaffffdfdaffff841affff841a000020260000202600007be6;
    assign coff[1685] = 256'h000040e0ffff91a9ffff91a9ffffbf20ffffbf2000006e5700006e57000040e0;
    assign coff[1686] = 256'h0000662affffb2e3ffffb2e3ffff99d6ffff99d600004d1d00004d1d0000662a;
    assign coff[1687] = 256'h000011b6ffff813bffff813bffffee4affffee4a00007ec500007ec5000011b6;
    assign coff[1688] = 256'h00007e74ffffec27ffffec27ffff818cffff818c000013d9000013d900007e74;
    assign coff[1689] = 256'h00004b61ffff988dffff988dffffb49fffffb49f000067730000677300004b61;
    assign coff[1690] = 256'h00006d3bffffbd45ffffbd45ffff92c5ffff92c5000042bb000042bb00006d3b;
    assign coff[1691] = 256'h00001e0effff8394ffff8394ffffe1f2ffffe1f200007c6c00007c6c00001e0e;
    assign coff[1692] = 256'h00007826ffffd3ddffffd3ddffff87daffff87da00002c2300002c2300007826;
    assign coff[1693] = 256'h000035c0ffff8bd5ffff8bd5ffffca40ffffca400000742b0000742b000035c0;
    assign coff[1694] = 256'h00005e1dffffa93effffa93effffa1e3ffffa1e3000056c2000056c200005e1d;
    assign coff[1695] = 256'h00000534ffff801bffff801bfffffaccfffffacc00007fe500007fe500000534;
    assign coff[1696] = 256'h00007feefffffbc7fffffbc7ffff8012ffff8012000004390000043900007fee;
    assign coff[1697] = 256'h0000577affffa28effffa28effffa886ffffa88600005d7200005d720000577a;
    assign coff[1698] = 256'h00007494ffffcb25ffffcb25ffff8b6cffff8b6c000034db000034db00007494;
    assign coff[1699] = 256'h00002d0fffff8831ffff8831ffffd2f1ffffd2f1000077cf000077cf00002d0f;
    assign coff[1700] = 256'h00007ca6ffffe2e7ffffe2e7ffff835affff835a00001d1900001d1900007ca6;
    assign coff[1701] = 256'h00004391ffff9349ffff9349ffffbc6fffffbc6f00006cb700006cb700004391;
    assign coff[1702] = 256'h00006806ffffb56bffffb56bffff97faffff97fa00004a9500004a9500006806;
    assign coff[1703] = 256'h000014d1ffff81b4ffff81b4ffffeb2fffffeb2f00007e4c00007e4c000014d1;
    assign coff[1704] = 256'h00007ee7ffffef43ffffef43ffff8119ffff8119000010bd000010bd00007ee7;
    assign coff[1705] = 256'h00004de5ffff9a6effff9a6effffb21bffffb21b000065920000659200004de5;
    assign coff[1706] = 256'h00006ed6ffffbff9ffffbff9ffff912affff912a000040070000400700006ed6;
    assign coff[1707] = 256'h00002119ffff845affff845affffdee7ffffdee700007ba600007ba600002119;
    assign coff[1708] = 256'h00007932ffffd6d3ffffd6d3ffff86ceffff86ce0000292d0000292d00007932;
    assign coff[1709] = 256'h00003895ffff8d30ffff8d30ffffc76bffffc76b000072d0000072d000003895;
    assign coff[1710] = 256'h00006037ffffab94ffffab94ffff9fc9ffff9fc90000546c0000546c00006037;
    assign coff[1711] = 256'h00000857ffff8046ffff8046fffff7a9fffff7a900007fba00007fba00000857;
    assign coff[1712] = 256'h00007f92fffff582fffff582ffff806effff806e00000a7e00000a7e00007f92;
    assign coff[1713] = 256'h000052c9ffff9e60ffff9e60ffffad37ffffad37000061a0000061a0000052c9;
    assign coff[1714] = 256'h000071d8ffffc57dffffc57dffff8e28ffff8e2800003a8300003a83000071d8;
    assign coff[1715] = 256'h00002720ffff8620ffff8620ffffd8e0ffffd8e0000079e0000079e000002720;
    assign coff[1716] = 256'h00007b12ffffdcd2ffffdcd2ffff84eeffff84ee0000232e0000232e00007b12;
    assign coff[1717] = 256'h00003e26ffff901affff901affffc1daffffc1da00006fe600006fe600003e26;
    assign coff[1718] = 256'h0000643effffb067ffffb067ffff9bc2ffff9bc200004f9900004f990000643e;
    assign coff[1719] = 256'h00000e99ffff80d6ffff80d6fffff167fffff16700007f2a00007f2a00000e99;
    assign coff[1720] = 256'h00007dedffffe90effffe90effff8213ffff8213000016f2000016f200007ded;
    assign coff[1721] = 256'h000048d1ffff96bbffff96bbffffb72fffffb72f0000694500006945000048d1;
    assign coff[1722] = 256'h00006b8fffffba9cffffba9cffff9471ffff9471000045640000456400006b8f;
    assign coff[1723] = 256'h00001afeffff82e1ffff82e1ffffe502ffffe50200007d1f00007d1f00001afe;
    assign coff[1724] = 256'h00007708ffffd0edffffd0edffff88f8ffff88f800002f1300002f1300007708;
    assign coff[1725] = 256'h000032e2ffff8a8cffff8a8cffffcd1effffcd1e0000757400007574000032e2;
    assign coff[1726] = 256'h00005bf5ffffa6f6ffffa6f6ffffa40bffffa40b0000590a0000590a00005bf5;
    assign coff[1727] = 256'h00000210ffff8004ffff8004fffffdf0fffffdf000007ffc00007ffc00000210;
    assign coff[1728] = 256'h00007ff9fffffd59fffffd59ffff8007ffff8007000002a7000002a700007ff9;
    assign coff[1729] = 256'h0000589effffa3a3ffffa3a3ffffa762ffffa76200005c5d00005c5d0000589e;
    assign coff[1730] = 256'h00007538ffffcc94ffffcc94ffff8ac8ffff8ac80000336c0000336c00007538;
    assign coff[1731] = 256'h00002e86ffff88c1ffff88c1ffffd17affffd17a0000773f0000773f00002e86;
    assign coff[1732] = 256'h00007cffffffe46fffffe46fffff8301ffff830100001b9100001b9100007cff;
    assign coff[1733] = 256'h000044e5ffff941fffff941fffffbb1bffffbb1b00006be100006be1000044e5;
    assign coff[1734] = 256'h000068efffffb6b3ffffb6b3ffff9711ffff97110000494d0000494d000068ef;
    assign coff[1735] = 256'h0000165effff81f8ffff81f8ffffe9a2ffffe9a200007e0800007e080000165e;
    assign coff[1736] = 256'h00007f19fffff0d2fffff0d2ffff80e7ffff80e700000f2e00000f2e00007f19;
    assign coff[1737] = 256'h00004f23ffff9b65ffff9b65ffffb0ddffffb0dd0000649b0000649b00004f23;
    assign coff[1738] = 256'h00006f9dffffc156ffffc156ffff9063ffff906300003eaa00003eaa00006f9d;
    assign coff[1739] = 256'h0000229dffff84c5ffff84c5ffffdd63ffffdd6300007b3b00007b3b0000229d;
    assign coff[1740] = 256'h000079b1ffffd851ffffd851ffff864fffff864f000027af000027af000079b1;
    assign coff[1741] = 256'h000039fdffff8de4ffff8de4ffffc603ffffc6030000721c0000721c000039fd;
    assign coff[1742] = 256'h0000613effffacc4ffffacc4ffff9ec2ffff9ec20000533c0000533c0000613e;
    assign coff[1743] = 256'h000009e8ffff8062ffff8062fffff618fffff61800007f9e00007f9e000009e8;
    assign coff[1744] = 256'h00007fb0fffff713fffff713ffff8050ffff8050000008ed000008ed00007fb0;
    assign coff[1745] = 256'h000053faffff9f66ffff9f66ffffac06ffffac060000609a0000609a000053fa;
    assign coff[1746] = 256'h0000728dffffc6e3ffffc6e3ffff8d73ffff8d730000391d0000391d0000728d;
    assign coff[1747] = 256'h0000289effff869effff869effffd762ffffd76200007962000079620000289e;
    assign coff[1748] = 256'h00007b7effffde56ffffde56ffff8482ffff8482000021aa000021aa00007b7e;
    assign coff[1749] = 256'h00003f85ffff90dfffff90dfffffc07bffffc07b00006f2100006f2100003f85;
    assign coff[1750] = 256'h00006536ffffb1a3ffffb1a3ffff9acaffff9aca00004e5d00004e5d00006536;
    assign coff[1751] = 256'h00001028ffff8106ffff8106ffffefd8ffffefd800007efa00007efa00001028;
    assign coff[1752] = 256'h00007e33ffffea9affffea9affff81cdffff81cd000015660000156600007e33;
    assign coff[1753] = 256'h00004a1bffff97a2ffff97a2ffffb5e5ffffb5e50000685e0000685e00004a1b;
    assign coff[1754] = 256'h00006c67ffffbbefffffbbefffff9399ffff9399000044110000441100006c67;
    assign coff[1755] = 256'h00001c86ffff8338ffff8338ffffe37affffe37a00007cc800007cc800001c86;
    assign coff[1756] = 256'h00007799ffffd264ffffd264ffff8867ffff886700002d9c00002d9c00007799;
    assign coff[1757] = 256'h00003452ffff8b2effff8b2effffcbaeffffcbae000074d2000074d200003452;
    assign coff[1758] = 256'h00005d0bffffa818ffffa818ffffa2f5ffffa2f5000057e8000057e800005d0b;
    assign coff[1759] = 256'h000003a2ffff800dffff800dfffffc5efffffc5e00007ff300007ff3000003a2;
    assign coff[1760] = 256'h00007fdefffffa36fffffa36ffff8022ffff8022000005ca000005ca00007fde;
    assign coff[1761] = 256'h00005653ffffa17dffffa17dffffa9adffffa9ad00005e8300005e8300005653;
    assign coff[1762] = 256'h000073ebffffc9b8ffffc9b8ffff8c15ffff8c150000364800003648000073eb;
    assign coff[1763] = 256'h00002b95ffff87a6ffff87a6ffffd46bffffd46b0000785a0000785a00002b95;
    assign coff[1764] = 256'h00007c48ffffe160ffffe160ffff83b8ffff83b800001ea000001ea000007c48;
    assign coff[1765] = 256'h0000423affff9277ffff9277ffffbdc6ffffbdc600006d8900006d890000423a;
    assign coff[1766] = 256'h0000671affffb425ffffb425ffff98e6ffff98e600004bdb00004bdb0000671a;
    assign coff[1767] = 256'h00001344ffff8175ffff8175ffffecbcffffecbc00007e8b00007e8b00001344;
    assign coff[1768] = 256'h00007eb0ffffedb4ffffedb4ffff8150ffff81500000124c0000124c00007eb0;
    assign coff[1769] = 256'h00004ca5ffff997cffff997cffffb35bffffb35b000066840000668400004ca5;
    assign coff[1770] = 256'h00006e0affffbe9effffbe9effff91f6ffff91f6000041620000416200006e0a;
    assign coff[1771] = 256'h00001f94ffff83f5ffff83f5ffffe06cffffe06c00007c0b00007c0b00001f94;
    assign coff[1772] = 256'h000078afffffd557ffffd557ffff8751ffff875100002aa900002aa9000078af;
    assign coff[1773] = 256'h0000372cffff8c80ffff8c80ffffc8d4ffffc8d400007380000073800000372c;
    assign coff[1774] = 256'h00005f2cffffaa68ffffaa68ffffa0d4ffffa0d4000055980000559800005f2c;
    assign coff[1775] = 256'h000006c5ffff802effff802efffff93bfffff93b00007fd200007fd2000006c5;
    assign coff[1776] = 256'h00007f6efffff3f1fffff3f1ffff8092ffff809200000c0f00000c0f00007f6e;
    assign coff[1777] = 256'h00005195ffff9d5effff9d5effffae6bffffae6b000062a2000062a200005195;
    assign coff[1778] = 256'h0000711effffc418ffffc418ffff8ee2ffff8ee200003be800003be80000711e;
    assign coff[1779] = 256'h000025a0ffff85a8ffff85a8ffffda60ffffda6000007a5800007a58000025a0;
    assign coff[1780] = 256'h00007aa1ffffdb50ffffdb50ffff855fffff855f000024b0000024b000007aa1;
    assign coff[1781] = 256'h00003cc5ffff8f59ffff8f59ffffc33bffffc33b000070a7000070a700003cc5;
    assign coff[1782] = 256'h00006342ffffaf2dffffaf2dffff9cbeffff9cbe000050d3000050d300006342;
    assign coff[1783] = 256'h00000d09ffff80aaffff80aafffff2f7fffff2f700007f5600007f5600000d09;
    assign coff[1784] = 256'h00007da3ffffe783ffffe783ffff825dffff825d0000187d0000187d00007da3;
    assign coff[1785] = 256'h00004785ffff95d8ffff95d8ffffb87bffffb87b00006a2800006a2800004785;
    assign coff[1786] = 256'h00006ab3ffffb94cffffb94cffff954dffff954d000046b4000046b400006ab3;
    assign coff[1787] = 256'h00001974ffff828effff828effffe68cffffe68c00007d7200007d7200001974;
    assign coff[1788] = 256'h00007672ffffcf78ffffcf78ffff898effff898e000030880000308800007672;
    assign coff[1789] = 256'h00003170ffff89efffff89efffffce90ffffce90000076110000761100003170;
    assign coff[1790] = 256'h00005adbffffa5d7ffffa5d7ffffa525ffffa52500005a2900005a2900005adb;
    assign coff[1791] = 256'h0000007effff8001ffff8001ffffff82ffffff8200007fff00007fff0000007e;
    assign coff[1792] = 256'h00007fffffffff50ffffff50ffff8001ffff8001000000b0000000b000007fff;
    assign coff[1793] = 256'h00005a06ffffa501ffffa501ffffa5faffffa5fa00005aff00005aff00005a06;
    assign coff[1794] = 256'h000075feffffce62ffffce62ffff8a02ffff8a020000319e0000319e000075fe;
    assign coff[1795] = 256'h00003059ffff897bffff897bffffcfa7ffffcfa7000076850000768500003059;
    assign coff[1796] = 256'h00007d68ffffe65bffffe65bffff8298ffff8298000019a5000019a500007d68;
    assign coff[1797] = 256'h0000468affff9531ffff9531ffffb976ffffb97600006acf00006acf0000468a;
    assign coff[1798] = 256'h00006a0bffffb851ffffb851ffff95f5ffff95f5000047af000047af00006a0b;
    assign coff[1799] = 256'h0000184cffff8254ffff8254ffffe7b4ffffe7b400007dac00007dac0000184c;
    assign coff[1800] = 256'h00007f50fffff2c5fffff2c5ffff80b0ffff80b000000d3b00000d3b00007f50;
    assign coff[1801] = 256'h000050acffff9c9fffff9c9fffffaf54ffffaf540000636100006361000050ac;
    assign coff[1802] = 256'h0000708fffffc30effffc30effff8f71ffff8f7100003cf200003cf20000708f;
    assign coff[1803] = 256'h00002480ffff8550ffff8550ffffdb80ffffdb8000007ab000007ab000002480;
    assign coff[1804] = 256'h00007a49ffffda30ffffda30ffff85b7ffff85b7000025d0000025d000007a49;
    assign coff[1805] = 256'h00003bbbffff8ecbffff8ecbffffc445ffffc445000071350000713500003bbb;
    assign coff[1806] = 256'h00006282ffffae45ffffae45ffff9d7effff9d7e000051bb000051bb00006282;
    assign coff[1807] = 256'h00000bddffff808dffff808dfffff423fffff42300007f7300007f7300000bdd;
    assign coff[1808] = 256'h00007fcffffff908fffff908ffff8031ffff8031000006f8000006f800007fcf;
    assign coff[1809] = 256'h00005573ffffa0b3ffffa0b3ffffaa8dffffaa8d00005f4d00005f4d00005573;
    assign coff[1810] = 256'h0000736affffc8a7ffffc8a7ffff8c96ffff8c9600003759000037590000736a;
    assign coff[1811] = 256'h00002a79ffff8741ffff8741ffffd587ffffd587000078bf000078bf00002a79;
    assign coff[1812] = 256'h00007bffffffe03bffffe03bffff8401ffff840100001fc500001fc500007bff;
    assign coff[1813] = 256'h00004137ffff91dcffff91dcffffbec9ffffbec900006e2400006e2400004137;
    assign coff[1814] = 256'h00006666ffffb333ffffb333ffff999affff999a00004ccd00004ccd00006666;
    assign coff[1815] = 256'h0000121affff8149ffff8149ffffede6ffffede600007eb700007eb70000121a;
    assign coff[1816] = 256'h00007e83ffffec8affffec8affff817dffff817d000013760000137600007e83;
    assign coff[1817] = 256'h00004bb2ffff98c8ffff98c8ffffb44effffb44e000067380000673800004bb2;
    assign coff[1818] = 256'h00006d6fffffbd9bffffbd9bffff9291ffff9291000042650000426500006d6f;
    assign coff[1819] = 256'h00001e6fffff83acffff83acffffe191ffffe19100007c5400007c5400001e6f;
    assign coff[1820] = 256'h00007849ffffd43bffffd43bffff87b7ffff87b700002bc500002bc500007849;
    assign coff[1821] = 256'h0000361bffff8bffffff8bffffffc9e5ffffc9e500007401000074010000361b;
    assign coff[1822] = 256'h00005e61ffffa988ffffa988ffffa19fffffa19f000056780000567800005e61;
    assign coff[1823] = 256'h00000598ffff801fffff801ffffffa68fffffa6800007fe100007fe100000598;
    assign coff[1824] = 256'h00007ff1fffffc2cfffffc2cffff800fffff800f000003d4000003d400007ff1;
    assign coff[1825] = 256'h000057c3ffffa2d3ffffa2d3ffffa83dffffa83d00005d2d00005d2d000057c3;
    assign coff[1826] = 256'h000074bdffffcb80ffffcb80ffff8b43ffff8b430000348000003480000074bd;
    assign coff[1827] = 256'h00002d6dffff8855ffff8855ffffd293ffffd293000077ab000077ab00002d6d;
    assign coff[1828] = 256'h00007cbdffffe349ffffe349ffff8343ffff834300001cb700001cb700007cbd;
    assign coff[1829] = 256'h000043e6ffff937effff937effffbc1affffbc1a00006c8200006c82000043e6;
    assign coff[1830] = 256'h00006841ffffb5bcffffb5bcffff97bfffff97bf00004a4400004a4400006841;
    assign coff[1831] = 256'h00001535ffff81c5ffff81c5ffffeacbffffeacb00007e3b00007e3b00001535;
    assign coff[1832] = 256'h00007ef4ffffefa6ffffefa6ffff810cffff810c0000105a0000105a00007ef4;
    assign coff[1833] = 256'h00004e35ffff9aacffff9aacffffb1cbffffb1cb000065540000655400004e35;
    assign coff[1834] = 256'h00006f08ffffc050ffffc050ffff90f8ffff90f800003fb000003fb000006f08;
    assign coff[1835] = 256'h0000217affff8475ffff8475ffffde86ffffde8600007b8b00007b8b0000217a;
    assign coff[1836] = 256'h00007953ffffd732ffffd732ffff86adffff86ad000028ce000028ce00007953;
    assign coff[1837] = 256'h000038f0ffff8d5cffff8d5cffffc710ffffc710000072a4000072a4000038f0;
    assign coff[1838] = 256'h00006079ffffabe0ffffabe0ffff9f87ffff9f87000054200000542000006079;
    assign coff[1839] = 256'h000008bbffff804cffff804cfffff745fffff74500007fb400007fb4000008bb;
    assign coff[1840] = 256'h00007f9afffff5e6fffff5e6ffff8066ffff806600000a1a00000a1a00007f9a;
    assign coff[1841] = 256'h00005316ffff9ea1ffff9ea1ffffaceaffffacea0000615f0000615f00005316;
    assign coff[1842] = 256'h00007206ffffc5d6ffffc5d6ffff8dfaffff8dfa00003a2a00003a2a00007206;
    assign coff[1843] = 256'h00002780ffff863fffff863fffffd880ffffd880000079c1000079c100002780;
    assign coff[1844] = 256'h00007b2effffdd33ffffdd33ffff84d2ffff84d2000022cd000022cd00007b2e;
    assign coff[1845] = 256'h00003e7effff904bffff904bffffc182ffffc18200006fb500006fb500003e7e;
    assign coff[1846] = 256'h0000647cffffb0b6ffffb0b6ffff9b84ffff9b8400004f4a00004f4a0000647c;
    assign coff[1847] = 256'h00000efcffff80e1ffff80e1fffff104fffff10400007f1f00007f1f00000efc;
    assign coff[1848] = 256'h00007dffffffe971ffffe971ffff8201ffff82010000168f0000168f00007dff;
    assign coff[1849] = 256'h00004924ffff96f4ffff96f4ffffb6dcffffb6dc0000690c0000690c00004924;
    assign coff[1850] = 256'h00006bc6ffffbaf1ffffbaf1ffff943affff943a0000450f0000450f00006bc6;
    assign coff[1851] = 256'h00001b60ffff82f6ffff82f6ffffe4a0ffffe4a000007d0a00007d0a00001b60;
    assign coff[1852] = 256'h0000772dffffd14bffffd14bffff88d3ffff88d300002eb500002eb50000772d;
    assign coff[1853] = 256'h0000333effff8ab4ffff8ab4ffffccc2ffffccc20000754c0000754c0000333e;
    assign coff[1854] = 256'h00005c3affffa73effffa73effffa3c6ffffa3c6000058c2000058c200005c3a;
    assign coff[1855] = 256'h00000274ffff8006ffff8006fffffd8cfffffd8c00007ffa00007ffa00000274;
    assign coff[1856] = 256'h00007ffbfffffdbefffffdbeffff8005ffff8005000002420000024200007ffb;
    assign coff[1857] = 256'h000058e6ffffa3e8ffffa3e8ffffa71affffa71a00005c1800005c18000058e6;
    assign coff[1858] = 256'h00007560ffffccf0ffffccf0ffff8aa0ffff8aa0000033100000331000007560;
    assign coff[1859] = 256'h00002ee4ffff88e6ffff88e6ffffd11cffffd11c0000771a0000771a00002ee4;
    assign coff[1860] = 256'h00007d15ffffe4d1ffffe4d1ffff82ebffff82eb00001b2f00001b2f00007d15;
    assign coff[1861] = 256'h00004539ffff9456ffff9456ffffbac7ffffbac700006baa00006baa00004539;
    assign coff[1862] = 256'h00006928ffffb705ffffb705ffff96d8ffff96d8000048fb000048fb00006928;
    assign coff[1863] = 256'h000016c1ffff820affff820affffe93fffffe93f00007df600007df6000016c1;
    assign coff[1864] = 256'h00007f24fffff135fffff135ffff80dcffff80dc00000ecb00000ecb00007f24;
    assign coff[1865] = 256'h00004f72ffff9ba3ffff9ba3ffffb08effffb08e0000645d0000645d00004f72;
    assign coff[1866] = 256'h00006fceffffc1aeffffc1aeffff9032ffff903200003e5200003e5200006fce;
    assign coff[1867] = 256'h000022fdffff84e0ffff84e0ffffdd03ffffdd0300007b2000007b20000022fd;
    assign coff[1868] = 256'h000079d0ffffd8b0ffffd8b0ffff8630ffff86300000275000002750000079d0;
    assign coff[1869] = 256'h00003a57ffff8e11ffff8e11ffffc5a9ffffc5a9000071ef000071ef00003a57;
    assign coff[1870] = 256'h0000617fffffad11ffffad11ffff9e81ffff9e81000052ef000052ef0000617f;
    assign coff[1871] = 256'h00000a4cffff806affff806afffff5b4fffff5b400007f9600007f9600000a4c;
    assign coff[1872] = 256'h00007fb7fffff777fffff777ffff8049ffff8049000008890000088900007fb7;
    assign coff[1873] = 256'h00005446ffff9fa8ffff9fa8ffffabbaffffabba000060580000605800005446;
    assign coff[1874] = 256'h000072baffffc73effffc73effff8d46ffff8d46000038c2000038c2000072ba;
    assign coff[1875] = 256'h000028fdffff86beffff86beffffd703ffffd7030000794200007942000028fd;
    assign coff[1876] = 256'h00007b99ffffdeb7ffffdeb7ffff8467ffff8467000021490000214900007b99;
    assign coff[1877] = 256'h00003fdcffff9111ffff9111ffffc024ffffc02400006eef00006eef00003fdc;
    assign coff[1878] = 256'h00006573ffffb1f3ffffb1f3ffff9a8dffff9a8d00004e0d00004e0d00006573;
    assign coff[1879] = 256'h0000108cffff8113ffff8113ffffef74ffffef7400007eed00007eed0000108c;
    assign coff[1880] = 256'h00007e43ffffeafdffffeafdffff81bdffff81bd000015030000150300007e43;
    assign coff[1881] = 256'h00004a6dffff97dcffff97dcffffb593ffffb593000068240000682400004a6d;
    assign coff[1882] = 256'h00006c9dffffbc45ffffbc45ffff9363ffff9363000043bb000043bb00006c9d;
    assign coff[1883] = 256'h00001ce8ffff834fffff834fffffe318ffffe31800007cb100007cb100001ce8;
    assign coff[1884] = 256'h000077bdffffd2c2ffffd2c2ffff8843ffff884300002d3e00002d3e000077bd;
    assign coff[1885] = 256'h000034adffff8b58ffff8b58ffffcb53ffffcb53000074a8000074a8000034ad;
    assign coff[1886] = 256'h00005d50ffffa861ffffa861ffffa2b0ffffa2b00000579f0000579f00005d50;
    assign coff[1887] = 256'h00000406ffff8010ffff8010fffffbfafffffbfa00007ff000007ff000000406;
    assign coff[1888] = 256'h00007fe3fffffa9afffffa9affff801dffff801d000005660000056600007fe3;
    assign coff[1889] = 256'h0000569dffffa1c1ffffa1c1ffffa963ffffa96300005e3f00005e3f0000569d;
    assign coff[1890] = 256'h00007416ffffca13ffffca13ffff8beaffff8bea000035ed000035ed00007416;
    assign coff[1891] = 256'h00002bf4ffff87c8ffff87c8ffffd40cffffd40c000078380000783800002bf4;
    assign coff[1892] = 256'h00007c60ffffe1c2ffffe1c2ffff83a0ffff83a000001e3e00001e3e00007c60;
    assign coff[1893] = 256'h00004290ffff92abffff92abffffbd70ffffbd7000006d5500006d5500004290;
    assign coff[1894] = 256'h00006756ffffb476ffffb476ffff98aaffff98aa00004b8a00004b8a00006756;
    assign coff[1895] = 256'h000013a8ffff8185ffff8185ffffec58ffffec5800007e7b00007e7b000013a8;
    assign coff[1896] = 256'h00007ebeffffee18ffffee18ffff8142ffff8142000011e8000011e800007ebe;
    assign coff[1897] = 256'h00004cf5ffff99b8ffff99b8ffffb30bffffb30b000066480000664800004cf5;
    assign coff[1898] = 256'h00006e3effffbef4ffffbef4ffff91c2ffff91c20000410c0000410c00006e3e;
    assign coff[1899] = 256'h00001ff5ffff840effff840effffe00bffffe00b00007bf200007bf200001ff5;
    assign coff[1900] = 256'h000078d0ffffd5b6ffffd5b6ffff8730ffff873000002a4a00002a4a000078d0;
    assign coff[1901] = 256'h00003786ffff8cabffff8cabffffc87affffc87a000073550000735500003786;
    assign coff[1902] = 256'h00005f6fffffaab2ffffaab2ffffa091ffffa0910000554e0000554e00005f6f;
    assign coff[1903] = 256'h0000072affff8033ffff8033fffff8d6fffff8d600007fcd00007fcd0000072a;
    assign coff[1904] = 256'h00007f78fffff455fffff455ffff8088ffff808800000bab00000bab00007f78;
    assign coff[1905] = 256'h000051e2ffff9d9effff9d9effffae1effffae1e0000626200006262000051e2;
    assign coff[1906] = 256'h0000714dffffc471ffffc471ffff8eb3ffff8eb300003b8f00003b8f0000714d;
    assign coff[1907] = 256'h00002600ffff85c5ffff85c5ffffda00ffffda0000007a3b00007a3b00002600;
    assign coff[1908] = 256'h00007abeffffdbb1ffffdbb1ffff8542ffff85420000244f0000244f00007abe;
    assign coff[1909] = 256'h00003d1effff8f89ffff8f89ffffc2e2ffffc2e2000070770000707700003d1e;
    assign coff[1910] = 256'h00006381ffffaf7cffffaf7cffff9c7fffff9c7f000050840000508400006381;
    assign coff[1911] = 256'h00000d6dffff80b5ffff80b5fffff293fffff29300007f4b00007f4b00000d6d;
    assign coff[1912] = 256'h00007db6ffffe7e5ffffe7e5ffff824affff824a0000181b0000181b00007db6;
    assign coff[1913] = 256'h000047d9ffff9611ffff9611ffffb827ffffb827000069ef000069ef000047d9;
    assign coff[1914] = 256'h00006aebffffb9a0ffffb9a0ffff9515ffff9515000046600000466000006aeb;
    assign coff[1915] = 256'h000019d6ffff82a3ffff82a3ffffe62affffe62a00007d5d00007d5d000019d6;
    assign coff[1916] = 256'h00007698ffffcfd6ffffcfd6ffff8968ffff89680000302a0000302a00007698;
    assign coff[1917] = 256'h000031ccffff8a16ffff8a16ffffce34ffffce34000075ea000075ea000031cc;
    assign coff[1918] = 256'h00005b22ffffa61effffa61effffa4deffffa4de000059e2000059e200005b22;
    assign coff[1919] = 256'h000000e2ffff8001ffff8001ffffff1effffff1e00007fff00007fff000000e2;
    assign coff[1920] = 256'h00007ffefffffe87fffffe87ffff8002ffff8002000001790000017900007ffe;
    assign coff[1921] = 256'h00005976ffffa474ffffa474ffffa68affffa68a00005b8c00005b8c00005976;
    assign coff[1922] = 256'h000075afffffcda9ffffcda9ffff8a51ffff8a510000325700003257000075af;
    assign coff[1923] = 256'h00002f9fffff8930ffff8930ffffd061ffffd061000076d0000076d000002f9f;
    assign coff[1924] = 256'h00007d3fffffe596ffffe596ffff82c1ffff82c100001a6a00001a6a00007d3f;
    assign coff[1925] = 256'h000045e2ffff94c3ffff94c3ffffba1effffba1e00006b3d00006b3d000045e2;
    assign coff[1926] = 256'h0000699affffb7abffffb7abffff9666ffff966600004855000048550000699a;
    assign coff[1927] = 256'h00001787ffff822effff822effffe879ffffe87900007dd200007dd200001787;
    assign coff[1928] = 256'h00007f3bfffff1fdfffff1fdffff80c5ffff80c500000e0300000e0300007f3b;
    assign coff[1929] = 256'h0000500fffff9c21ffff9c21ffffaff1ffffaff1000063df000063df0000500f;
    assign coff[1930] = 256'h0000702fffffc25effffc25effff8fd1ffff8fd100003da200003da20000702f;
    assign coff[1931] = 256'h000023bfffff8518ffff8518ffffdc41ffffdc4100007ae800007ae8000023bf;
    assign coff[1932] = 256'h00007a0effffd970ffffd970ffff85f2ffff85f2000026900000269000007a0e;
    assign coff[1933] = 256'h00003b09ffff8e6dffff8e6dffffc4f7ffffc4f7000071930000719300003b09;
    assign coff[1934] = 256'h00006201ffffadaaffffadaaffff9dffffff9dff000052560000525600006201;
    assign coff[1935] = 256'h00000b14ffff807bffff807bfffff4ecfffff4ec00007f8500007f8500000b14;
    assign coff[1936] = 256'h00007fc4fffff840fffff840ffff803cffff803c000007c0000007c000007fc4;
    assign coff[1937] = 256'h000054ddffffa02dffffa02dffffab23ffffab2300005fd300005fd3000054dd;
    assign coff[1938] = 256'h00007313ffffc7f2ffffc7f2ffff8cedffff8ced0000380e0000380e00007313;
    assign coff[1939] = 256'h000029bcffff86ffffff86ffffffd644ffffd6440000790100007901000029bc;
    assign coff[1940] = 256'h00007bccffffdf79ffffdf79ffff8434ffff8434000020870000208700007bcc;
    assign coff[1941] = 256'h0000408affff9176ffff9176ffffbf76ffffbf7600006e8a00006e8a0000408a;
    assign coff[1942] = 256'h000065edffffb293ffffb293ffff9a13ffff9a1300004d6d00004d6d000065ed;
    assign coff[1943] = 256'h00001153ffff812dffff812dffffeeadffffeead00007ed300007ed300001153;
    assign coff[1944] = 256'h00007e64ffffebc3ffffebc3ffff819cffff819c0000143d0000143d00007e64;
    assign coff[1945] = 256'h00004b10ffff9852ffff9852ffffb4f0ffffb4f0000067ae000067ae00004b10;
    assign coff[1946] = 256'h00006d06ffffbcf0ffffbcf0ffff92faffff92fa000043100000431000006d06;
    assign coff[1947] = 256'h00001dacffff837dffff837dffffe254ffffe25400007c8300007c8300001dac;
    assign coff[1948] = 256'h00007803ffffd37fffffd37fffff87fdffff87fd00002c8100002c8100007803;
    assign coff[1949] = 256'h00003564ffff8babffff8babffffca9cffffca9c000074550000745500003564;
    assign coff[1950] = 256'h00005dd9ffffa8f4ffffa8f4ffffa227ffffa2270000570c0000570c00005dd9;
    assign coff[1951] = 256'h000004cfffff8017ffff8017fffffb31fffffb3100007fe900007fe9000004cf;
    assign coff[1952] = 256'h00007febfffffb63fffffb63ffff8015ffff80150000049d0000049d00007feb;
    assign coff[1953] = 256'h00005730ffffa249ffffa249ffffa8d0ffffa8d000005db700005db700005730;
    assign coff[1954] = 256'h0000746affffcac9ffffcac9ffff8b96ffff8b9600003537000035370000746a;
    assign coff[1955] = 256'h00002cb1ffff880effff880effffd34fffffd34f000077f2000077f200002cb1;
    assign coff[1956] = 256'h00007c8fffffe285ffffe285ffff8371ffff837100001d7b00001d7b00007c8f;
    assign coff[1957] = 256'h0000433bffff9314ffff9314ffffbcc5ffffbcc500006cec00006cec0000433b;
    assign coff[1958] = 256'h000067ccffffb519ffffb519ffff9834ffff983400004ae700004ae7000067cc;
    assign coff[1959] = 256'h0000146effff81a4ffff81a4ffffeb92ffffeb9200007e5c00007e5c0000146e;
    assign coff[1960] = 256'h00007ed9ffffeedfffffeedfffff8127ffff8127000011210000112100007ed9;
    assign coff[1961] = 256'h00004d95ffff9a31ffff9a31ffffb26bffffb26b000065cf000065cf00004d95;
    assign coff[1962] = 256'h00006ea3ffffbfa2ffffbfa2ffff915dffff915d0000405e0000405e00006ea3;
    assign coff[1963] = 256'h000020b8ffff8441ffff8441ffffdf48ffffdf4800007bbf00007bbf000020b8;
    assign coff[1964] = 256'h00007912ffffd674ffffd674ffff86eeffff86ee0000298c0000298c00007912;
    assign coff[1965] = 256'h0000383bffff8d03ffff8d03ffffc7c5ffffc7c5000072fd000072fd0000383b;
    assign coff[1966] = 256'h00005ff4ffffab49ffffab49ffffa00cffffa00c000054b7000054b700005ff4;
    assign coff[1967] = 256'h000007f2ffff803fffff803ffffff80efffff80e00007fc100007fc1000007f2;
    assign coff[1968] = 256'h00007f89fffff51efffff51effff8077ffff807700000ae200000ae200007f89;
    assign coff[1969] = 256'h0000527cffff9e1fffff9e1fffffad84ffffad84000061e1000061e10000527c;
    assign coff[1970] = 256'h000071aaffffc523ffffc523ffff8e56ffff8e5600003add00003add000071aa;
    assign coff[1971] = 256'h000026c0ffff8602ffff8602ffffd940ffffd940000079fe000079fe000026c0;
    assign coff[1972] = 256'h00007af6ffffdc72ffffdc72ffff850affff850a0000238e0000238e00007af6;
    assign coff[1973] = 256'h00003dceffff8fe9ffff8fe9ffffc232ffffc232000070170000701700003dce;
    assign coff[1974] = 256'h000063ffffffb018ffffb018ffff9c01ffff9c0100004fe800004fe8000063ff;
    assign coff[1975] = 256'h00000e35ffff80caffff80cafffff1cbfffff1cb00007f3600007f3600000e35;
    assign coff[1976] = 256'h00007ddbffffe8abffffe8abffff8225ffff8225000017550000175500007ddb;
    assign coff[1977] = 256'h0000487fffff9682ffff9682ffffb781ffffb7810000697e0000697e0000487f;
    assign coff[1978] = 256'h00006b59ffffba48ffffba48ffff94a7ffff94a7000045b8000045b800006b59;
    assign coff[1979] = 256'h00001a9bffff82ccffff82ccffffe565ffffe56500007d3400007d3400001a9b;
    assign coff[1980] = 256'h000076e3ffffd090ffffd090ffff891dffff891d00002f7000002f70000076e3;
    assign coff[1981] = 256'h00003285ffff8a64ffff8a64ffffcd7bffffcd7b0000759c0000759c00003285;
    assign coff[1982] = 256'h00005bafffffa6aeffffa6aeffffa451ffffa451000059520000595200005baf;
    assign coff[1983] = 256'h000001abffff8003ffff8003fffffe55fffffe5500007ffd00007ffd000001ab;
    assign coff[1984] = 256'h00007ff7fffffcf5fffffcf5ffff8009ffff80090000030b0000030b00007ff7;
    assign coff[1985] = 256'h00005855ffffa35dffffa35dffffa7abffffa7ab00005ca300005ca300005855;
    assign coff[1986] = 256'h0000750fffffcc38ffffcc38ffff8af1ffff8af1000033c8000033c80000750f;
    assign coff[1987] = 256'h00002e28ffff889dffff889dffffd1d8ffffd1d8000077630000776300002e28;
    assign coff[1988] = 256'h00007ce9ffffe40dffffe40dffff8317ffff831700001bf300001bf300007ce9;
    assign coff[1989] = 256'h00004490ffff93e9ffff93e9ffffbb70ffffbb7000006c1700006c1700004490;
    assign coff[1990] = 256'h000068b5ffffb660ffffb660ffff974bffff974b000049a0000049a0000068b5;
    assign coff[1991] = 256'h000015fbffff81e7ffff81e7ffffea05ffffea0500007e1900007e19000015fb;
    assign coff[1992] = 256'h00007f0dfffff06efffff06effff80f3ffff80f300000f9200000f9200007f0d;
    assign coff[1993] = 256'h00004ed4ffff9b27ffff9b27ffffb12cffffb12c000064d9000064d900004ed4;
    assign coff[1994] = 256'h00006f6bffffc0ffffffc0ffffff9095ffff909500003f0100003f0100006f6b;
    assign coff[1995] = 256'h0000223cffff84aaffff84aaffffddc4ffffddc400007b5600007b560000223c;
    assign coff[1996] = 256'h00007992ffffd7f1ffffd7f1ffff866effff866e0000280f0000280f00007992;
    assign coff[1997] = 256'h000039a3ffff8db6ffff8db6ffffc65dffffc65d0000724a0000724a000039a3;
    assign coff[1998] = 256'h000060fdffffac78ffffac78ffff9f03ffff9f030000538800005388000060fd;
    assign coff[1999] = 256'h00000984ffff805bffff805bfffff67cfffff67c00007fa500007fa500000984;
    assign coff[2000] = 256'h00007fa9fffff6affffff6afffff8057ffff8057000009510000095100007fa9;
    assign coff[2001] = 256'h000053aeffff9f24ffff9f24ffffac52ffffac52000060dc000060dc000053ae;
    assign coff[2002] = 256'h00007260ffffc68affffc68affff8da0ffff8da0000039760000397600007260;
    assign coff[2003] = 256'h0000283fffff867effff867effffd7c1ffffd7c100007982000079820000283f;
    assign coff[2004] = 256'h00007b64ffffddf5ffffddf5ffff849cffff849c0000220b0000220b00007b64;
    assign coff[2005] = 256'h00003f2dffff90adffff90adffffc0d3ffffc0d300006f5300006f5300003f2d;
    assign coff[2006] = 256'h000064f8ffffb154ffffb154ffff9b08ffff9b0800004eac00004eac000064f8;
    assign coff[2007] = 256'h00000fc4ffff80faffff80fafffff03cfffff03c00007f0600007f0600000fc4;
    assign coff[2008] = 256'h00007e22ffffea37ffffea37ffff81deffff81de000015c9000015c900007e22;
    assign coff[2009] = 256'h000049c9ffff9768ffff9768ffffb637ffffb6370000689800006898000049c9;
    assign coff[2010] = 256'h00006c32ffffbb9affffbb9affff93ceffff93ce000044660000446600006c32;
    assign coff[2011] = 256'h00001c24ffff8322ffff8322ffffe3dcffffe3dc00007cde00007cde00001c24;
    assign coff[2012] = 256'h00007775ffffd206ffffd206ffff888bffff888b00002dfa00002dfa00007775;
    assign coff[2013] = 256'h000033f6ffff8b05ffff8b05ffffcc0affffcc0a000074fb000074fb000033f6;
    assign coff[2014] = 256'h00005cc5ffffa7cfffffa7cfffffa33bffffa33b000058310000583100005cc5;
    assign coff[2015] = 256'h0000033dffff800affff800afffffcc3fffffcc300007ff600007ff60000033d;
    assign coff[2016] = 256'h00007fdafffff9d1fffff9d1ffff8026ffff80260000062f0000062f00007fda;
    assign coff[2017] = 256'h00005608ffffa139ffffa139ffffa9f8ffffa9f800005ec700005ec700005608;
    assign coff[2018] = 256'h000073c1ffffc95dffffc95dffff8c3fffff8c3f000036a3000036a3000073c1;
    assign coff[2019] = 256'h00002b37ffff8784ffff8784ffffd4c9ffffd4c90000787c0000787c00002b37;
    assign coff[2020] = 256'h00007c30ffffe0feffffe0feffff83d0ffff83d000001f0200001f0200007c30;
    assign coff[2021] = 256'h000041e4ffff9243ffff9243ffffbe1cffffbe1c00006dbd00006dbd000041e4;
    assign coff[2022] = 256'h000066deffffb3d4ffffb3d4ffff9922ffff992200004c2c00004c2c000066de;
    assign coff[2023] = 256'h000012e1ffff8166ffff8166ffffed1fffffed1f00007e9a00007e9a000012e1;
    assign coff[2024] = 256'h00007ea1ffffed51ffffed51ffff815fffff815f000012af000012af00007ea1;
    assign coff[2025] = 256'h00004c54ffff993fffff993fffffb3acffffb3ac000066c1000066c100004c54;
    assign coff[2026] = 256'h00006dd7ffffbe47ffffbe47ffff9229ffff9229000041b9000041b900006dd7;
    assign coff[2027] = 256'h00001f32ffff83dcffff83dcffffe0ceffffe0ce00007c2400007c2400001f32;
    assign coff[2028] = 256'h0000788dffffd4f8ffffd4f8ffff8773ffff877300002b0800002b080000788d;
    assign coff[2029] = 256'h000036d1ffff8c55ffff8c55ffffc92fffffc92f000073ab000073ab000036d1;
    assign coff[2030] = 256'h00005ee8ffffaa1dffffaa1dffffa118ffffa118000055e3000055e300005ee8;
    assign coff[2031] = 256'h00000661ffff8029ffff8029fffff99ffffff99f00007fd700007fd700000661;
    assign coff[2032] = 256'h00007f65fffff38dfffff38dffff809bffff809b00000c7300000c7300007f65;
    assign coff[2033] = 256'h00005147ffff9d1effff9d1effffaeb9ffffaeb9000062e2000062e200005147;
    assign coff[2034] = 256'h000070efffffc3bfffffc3bfffff8f11ffff8f1100003c4100003c41000070ef;
    assign coff[2035] = 256'h00002540ffff858affff858affffdac0ffffdac000007a7600007a7600002540;
    assign coff[2036] = 256'h00007a84ffffdaf0ffffdaf0ffff857cffff857c000025100000251000007a84;
    assign coff[2037] = 256'h00003c6dffff8f29ffff8f29ffffc393ffffc393000070d7000070d700003c6d;
    assign coff[2038] = 256'h00006302ffffaee0ffffaee0ffff9cfeffff9cfe000051200000512000006302;
    assign coff[2039] = 256'h00000ca5ffff80a0ffff80a0fffff35bfffff35b00007f6000007f6000000ca5;
    assign coff[2040] = 256'h00007d8fffffe720ffffe720ffff8271ffff8271000018e0000018e000007d8f;
    assign coff[2041] = 256'h00004732ffff95a0ffff95a0ffffb8ceffffb8ce00006a6000006a6000004732;
    assign coff[2042] = 256'h00006a7cffffb8f8ffffb8f8ffff9584ffff9584000047080000470800006a7c;
    assign coff[2043] = 256'h00001911ffff827bffff827bffffe6efffffe6ef00007d8500007d8500001911;
    assign coff[2044] = 256'h0000764bffffcf1bffffcf1bffff89b5ffff89b5000030e5000030e50000764b;
    assign coff[2045] = 256'h00003113ffff89c8ffff89c8ffffceedffffceed000076380000763800003113;
    assign coff[2046] = 256'h00005a94ffffa58fffffa58fffffa56cffffa56c00005a7100005a7100005a94;
    assign coff[2047] = 256'h00000019ffff8001ffff8001ffffffe7ffffffe700007fff00007fff00000019;




    always_ff @(posedge clk, negedge rst_n) begin
        if(~rst_n) begin
            data_o <= 'b0;
        end else if (valid == 1) begin
            data_o <= coff[addr_i];
        end else begin
            data_o <= 'b0;
        end
    end


endmodule