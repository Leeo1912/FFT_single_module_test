`timescale 1ns/1ps
module rom_1_rfft_data64
(
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic                     valid,
    input  logic [10:0]              addr_col1,
    input  logic [10:0]              addr_col2,
    output logic [63:0]              data_o_col1,
    output logic [63:0]              data_o_col2
);

    logic [63:0] coff[2047:0];

    assign coff[0   ] = 64'h00007fff00000000;
    assign coff[1   ] = 64'h00007ffffffffff3;
    assign coff[2   ] = 64'h00007fffffffffe7;
    assign coff[3   ] = 64'h00007fffffffffda;
    assign coff[4   ] = 64'h00007fffffffffce;
    assign coff[5   ] = 64'h00007fffffffffc1;
    assign coff[6   ] = 64'h00007fffffffffb5;
    assign coff[7   ] = 64'h00007fffffffffa8;
    assign coff[8   ] = 64'h00007fffffffff9b;
    assign coff[9   ] = 64'h00007fffffffff8f;
    assign coff[10  ] = 64'h00007fffffffff82;
    assign coff[11  ] = 64'h00007fffffffff76;
    assign coff[12  ] = 64'h00007fffffffff69;
    assign coff[13  ] = 64'h00007fffffffff5d;
    assign coff[14  ] = 64'h00007fffffffff50;
    assign coff[15  ] = 64'h00007fffffffff44;
    assign coff[16  ] = 64'h00007fffffffff37;
    assign coff[17  ] = 64'h00007fffffffff2a;
    assign coff[18  ] = 64'h00007fffffffff1e;
    assign coff[19  ] = 64'h00007fffffffff11;
    assign coff[20  ] = 64'h00007fffffffff05;
    assign coff[21  ] = 64'h00007ffffffffef8;
    assign coff[22  ] = 64'h00007ffffffffeec;
    assign coff[23  ] = 64'h00007ffffffffedf;
    assign coff[24  ] = 64'h00007ffffffffed2;
    assign coff[25  ] = 64'h00007ffefffffec6;
    assign coff[26  ] = 64'h00007ffefffffeb9;
    assign coff[27  ] = 64'h00007ffefffffead;
    assign coff[28  ] = 64'h00007ffefffffea0;
    assign coff[29  ] = 64'h00007ffefffffe94;
    assign coff[30  ] = 64'h00007ffefffffe87;
    assign coff[31  ] = 64'h00007ffefffffe7a;
    assign coff[32  ] = 64'h00007ffefffffe6e;
    assign coff[33  ] = 64'h00007ffdfffffe61;
    assign coff[34  ] = 64'h00007ffdfffffe55;
    assign coff[35  ] = 64'h00007ffdfffffe48;
    assign coff[36  ] = 64'h00007ffdfffffe3c;
    assign coff[37  ] = 64'h00007ffdfffffe2f;
    assign coff[38  ] = 64'h00007ffdfffffe22;
    assign coff[39  ] = 64'h00007ffcfffffe16;
    assign coff[40  ] = 64'h00007ffcfffffe09;
    assign coff[41  ] = 64'h00007ffcfffffdfd;
    assign coff[42  ] = 64'h00007ffcfffffdf0;
    assign coff[43  ] = 64'h00007ffcfffffde4;
    assign coff[44  ] = 64'h00007ffbfffffdd7;
    assign coff[45  ] = 64'h00007ffbfffffdcb;
    assign coff[46  ] = 64'h00007ffbfffffdbe;
    assign coff[47  ] = 64'h00007ffbfffffdb1;
    assign coff[48  ] = 64'h00007ffafffffda5;
    assign coff[49  ] = 64'h00007ffafffffd98;
    assign coff[50  ] = 64'h00007ffafffffd8c;
    assign coff[51  ] = 64'h00007ffafffffd7f;
    assign coff[52  ] = 64'h00007ff9fffffd73;
    assign coff[53  ] = 64'h00007ff9fffffd66;
    assign coff[54  ] = 64'h00007ff9fffffd59;
    assign coff[55  ] = 64'h00007ff9fffffd4d;
    assign coff[56  ] = 64'h00007ff8fffffd40;
    assign coff[57  ] = 64'h00007ff8fffffd34;
    assign coff[58  ] = 64'h00007ff8fffffd27;
    assign coff[59  ] = 64'h00007ff8fffffd1b;
    assign coff[60  ] = 64'h00007ff7fffffd0e;
    assign coff[61  ] = 64'h00007ff7fffffd02;
    assign coff[62  ] = 64'h00007ff7fffffcf5;
    assign coff[63  ] = 64'h00007ff6fffffce8;
    assign coff[64  ] = 64'h00007ff6fffffcdc;
    assign coff[65  ] = 64'h00007ff6fffffccf;
    assign coff[66  ] = 64'h00007ff6fffffcc3;
    assign coff[67  ] = 64'h00007ff5fffffcb6;
    assign coff[68  ] = 64'h00007ff5fffffcaa;
    assign coff[69  ] = 64'h00007ff5fffffc9d;
    assign coff[70  ] = 64'h00007ff4fffffc90;
    assign coff[71  ] = 64'h00007ff4fffffc84;
    assign coff[72  ] = 64'h00007ff4fffffc77;
    assign coff[73  ] = 64'h00007ff3fffffc6b;
    assign coff[74  ] = 64'h00007ff3fffffc5e;
    assign coff[75  ] = 64'h00007ff2fffffc52;
    assign coff[76  ] = 64'h00007ff2fffffc45;
    assign coff[77  ] = 64'h00007ff2fffffc39;
    assign coff[78  ] = 64'h00007ff1fffffc2c;
    assign coff[79  ] = 64'h00007ff1fffffc1f;
    assign coff[80  ] = 64'h00007ff1fffffc13;
    assign coff[81  ] = 64'h00007ff0fffffc06;
    assign coff[82  ] = 64'h00007ff0fffffbfa;
    assign coff[83  ] = 64'h00007feffffffbed;
    assign coff[84  ] = 64'h00007feffffffbe1;
    assign coff[85  ] = 64'h00007feffffffbd4;
    assign coff[86  ] = 64'h00007feefffffbc7;
    assign coff[87  ] = 64'h00007feefffffbbb;
    assign coff[88  ] = 64'h00007fedfffffbae;
    assign coff[89  ] = 64'h00007fedfffffba2;
    assign coff[90  ] = 64'h00007fecfffffb95;
    assign coff[91  ] = 64'h00007fecfffffb89;
    assign coff[92  ] = 64'h00007fecfffffb7c;
    assign coff[93  ] = 64'h00007febfffffb70;
    assign coff[94  ] = 64'h00007febfffffb63;
    assign coff[95  ] = 64'h00007feafffffb56;
    assign coff[96  ] = 64'h00007feafffffb4a;
    assign coff[97  ] = 64'h00007fe9fffffb3d;
    assign coff[98  ] = 64'h00007fe9fffffb31;
    assign coff[99  ] = 64'h00007fe8fffffb24;
    assign coff[100 ] = 64'h00007fe8fffffb18;
    assign coff[101 ] = 64'h00007fe7fffffb0b;
    assign coff[102 ] = 64'h00007fe7fffffaff;
    assign coff[103 ] = 64'h00007fe6fffffaf2;
    assign coff[104 ] = 64'h00007fe6fffffae5;
    assign coff[105 ] = 64'h00007fe5fffffad9;
    assign coff[106 ] = 64'h00007fe5fffffacc;
    assign coff[107 ] = 64'h00007fe4fffffac0;
    assign coff[108 ] = 64'h00007fe4fffffab3;
    assign coff[109 ] = 64'h00007fe3fffffaa7;
    assign coff[110 ] = 64'h00007fe3fffffa9a;
    assign coff[111 ] = 64'h00007fe2fffffa8e;
    assign coff[112 ] = 64'h00007fe2fffffa81;
    assign coff[113 ] = 64'h00007fe1fffffa74;
    assign coff[114 ] = 64'h00007fe1fffffa68;
    assign coff[115 ] = 64'h00007fe0fffffa5b;
    assign coff[116 ] = 64'h00007fe0fffffa4f;
    assign coff[117 ] = 64'h00007fdffffffa42;
    assign coff[118 ] = 64'h00007fdefffffa36;
    assign coff[119 ] = 64'h00007fdefffffa29;
    assign coff[120 ] = 64'h00007fddfffffa1d;
    assign coff[121 ] = 64'h00007fddfffffa10;
    assign coff[122 ] = 64'h00007fdcfffffa03;
    assign coff[123 ] = 64'h00007fdcfffff9f7;
    assign coff[124 ] = 64'h00007fdbfffff9ea;
    assign coff[125 ] = 64'h00007fdafffff9de;
    assign coff[126 ] = 64'h00007fdafffff9d1;
    assign coff[127 ] = 64'h00007fd9fffff9c5;
    assign coff[128 ] = 64'h00007fd9fffff9b8;
    assign coff[129 ] = 64'h00007fd8fffff9ac;
    assign coff[130 ] = 64'h00007fd7fffff99f;
    assign coff[131 ] = 64'h00007fd7fffff992;
    assign coff[132 ] = 64'h00007fd6fffff986;
    assign coff[133 ] = 64'h00007fd5fffff979;
    assign coff[134 ] = 64'h00007fd5fffff96d;
    assign coff[135 ] = 64'h00007fd4fffff960;
    assign coff[136 ] = 64'h00007fd3fffff954;
    assign coff[137 ] = 64'h00007fd3fffff947;
    assign coff[138 ] = 64'h00007fd2fffff93b;
    assign coff[139 ] = 64'h00007fd1fffff92e;
    assign coff[140 ] = 64'h00007fd1fffff922;
    assign coff[141 ] = 64'h00007fd0fffff915;
    assign coff[142 ] = 64'h00007fcffffff908;
    assign coff[143 ] = 64'h00007fcffffff8fc;
    assign coff[144 ] = 64'h00007fcefffff8ef;
    assign coff[145 ] = 64'h00007fcdfffff8e3;
    assign coff[146 ] = 64'h00007fcdfffff8d6;
    assign coff[147 ] = 64'h00007fccfffff8ca;
    assign coff[148 ] = 64'h00007fcbfffff8bd;
    assign coff[149 ] = 64'h00007fcbfffff8b1;
    assign coff[150 ] = 64'h00007fcafffff8a4;
    assign coff[151 ] = 64'h00007fc9fffff898;
    assign coff[152 ] = 64'h00007fc8fffff88b;
    assign coff[153 ] = 64'h00007fc8fffff87e;
    assign coff[154 ] = 64'h00007fc7fffff872;
    assign coff[155 ] = 64'h00007fc6fffff865;
    assign coff[156 ] = 64'h00007fc5fffff859;
    assign coff[157 ] = 64'h00007fc5fffff84c;
    assign coff[158 ] = 64'h00007fc4fffff840;
    assign coff[159 ] = 64'h00007fc3fffff833;
    assign coff[160 ] = 64'h00007fc2fffff827;
    assign coff[161 ] = 64'h00007fc2fffff81a;
    assign coff[162 ] = 64'h00007fc1fffff80e;
    assign coff[163 ] = 64'h00007fc0fffff801;
    assign coff[164 ] = 64'h00007fbffffff7f4;
    assign coff[165 ] = 64'h00007fbefffff7e8;
    assign coff[166 ] = 64'h00007fbefffff7db;
    assign coff[167 ] = 64'h00007fbdfffff7cf;
    assign coff[168 ] = 64'h00007fbcfffff7c2;
    assign coff[169 ] = 64'h00007fbbfffff7b6;
    assign coff[170 ] = 64'h00007fbafffff7a9;
    assign coff[171 ] = 64'h00007fbafffff79d;
    assign coff[172 ] = 64'h00007fb9fffff790;
    assign coff[173 ] = 64'h00007fb8fffff784;
    assign coff[174 ] = 64'h00007fb7fffff777;
    assign coff[175 ] = 64'h00007fb6fffff76b;
    assign coff[176 ] = 64'h00007fb5fffff75e;
    assign coff[177 ] = 64'h00007fb5fffff751;
    assign coff[178 ] = 64'h00007fb4fffff745;
    assign coff[179 ] = 64'h00007fb3fffff738;
    assign coff[180 ] = 64'h00007fb2fffff72c;
    assign coff[181 ] = 64'h00007fb1fffff71f;
    assign coff[182 ] = 64'h00007fb0fffff713;
    assign coff[183 ] = 64'h00007faffffff706;
    assign coff[184 ] = 64'h00007faefffff6fa;
    assign coff[185 ] = 64'h00007faefffff6ed;
    assign coff[186 ] = 64'h00007fadfffff6e1;
    assign coff[187 ] = 64'h00007facfffff6d4;
    assign coff[188 ] = 64'h00007fabfffff6c8;
    assign coff[189 ] = 64'h00007faafffff6bb;
    assign coff[190 ] = 64'h00007fa9fffff6af;
    assign coff[191 ] = 64'h00007fa8fffff6a2;
    assign coff[192 ] = 64'h00007fa7fffff695;
    assign coff[193 ] = 64'h00007fa6fffff689;
    assign coff[194 ] = 64'h00007fa5fffff67c;
    assign coff[195 ] = 64'h00007fa4fffff670;
    assign coff[196 ] = 64'h00007fa3fffff663;
    assign coff[197 ] = 64'h00007fa3fffff657;
    assign coff[198 ] = 64'h00007fa2fffff64a;
    assign coff[199 ] = 64'h00007fa1fffff63e;
    assign coff[200 ] = 64'h00007fa0fffff631;
    assign coff[201 ] = 64'h00007f9ffffff625;
    assign coff[202 ] = 64'h00007f9efffff618;
    assign coff[203 ] = 64'h00007f9dfffff60c;
    assign coff[204 ] = 64'h00007f9cfffff5ff;
    assign coff[205 ] = 64'h00007f9bfffff5f3;
    assign coff[206 ] = 64'h00007f9afffff5e6;
    assign coff[207 ] = 64'h00007f99fffff5d9;
    assign coff[208 ] = 64'h00007f98fffff5cd;
    assign coff[209 ] = 64'h00007f97fffff5c0;
    assign coff[210 ] = 64'h00007f96fffff5b4;
    assign coff[211 ] = 64'h00007f95fffff5a7;
    assign coff[212 ] = 64'h00007f94fffff59b;
    assign coff[213 ] = 64'h00007f93fffff58e;
    assign coff[214 ] = 64'h00007f92fffff582;
    assign coff[215 ] = 64'h00007f91fffff575;
    assign coff[216 ] = 64'h00007f90fffff569;
    assign coff[217 ] = 64'h00007f8ffffff55c;
    assign coff[218 ] = 64'h00007f8efffff550;
    assign coff[219 ] = 64'h00007f8dfffff543;
    assign coff[220 ] = 64'h00007f8bfffff537;
    assign coff[221 ] = 64'h00007f8afffff52a;
    assign coff[222 ] = 64'h00007f89fffff51e;
    assign coff[223 ] = 64'h00007f88fffff511;
    assign coff[224 ] = 64'h00007f87fffff505;
    assign coff[225 ] = 64'h00007f86fffff4f8;
    assign coff[226 ] = 64'h00007f85fffff4ec;
    assign coff[227 ] = 64'h00007f84fffff4df;
    assign coff[228 ] = 64'h00007f83fffff4d3;
    assign coff[229 ] = 64'h00007f82fffff4c6;
    assign coff[230 ] = 64'h00007f81fffff4b9;
    assign coff[231 ] = 64'h00007f80fffff4ad;
    assign coff[232 ] = 64'h00007f7efffff4a0;
    assign coff[233 ] = 64'h00007f7dfffff494;
    assign coff[234 ] = 64'h00007f7cfffff487;
    assign coff[235 ] = 64'h00007f7bfffff47b;
    assign coff[236 ] = 64'h00007f7afffff46e;
    assign coff[237 ] = 64'h00007f79fffff462;
    assign coff[238 ] = 64'h00007f78fffff455;
    assign coff[239 ] = 64'h00007f76fffff449;
    assign coff[240 ] = 64'h00007f75fffff43c;
    assign coff[241 ] = 64'h00007f74fffff430;
    assign coff[242 ] = 64'h00007f73fffff423;
    assign coff[243 ] = 64'h00007f72fffff417;
    assign coff[244 ] = 64'h00007f71fffff40a;
    assign coff[245 ] = 64'h00007f6ffffff3fe;
    assign coff[246 ] = 64'h00007f6efffff3f1;
    assign coff[247 ] = 64'h00007f6dfffff3e5;
    assign coff[248 ] = 64'h00007f6cfffff3d8;
    assign coff[249 ] = 64'h00007f6bfffff3cc;
    assign coff[250 ] = 64'h00007f6afffff3bf;
    assign coff[251 ] = 64'h00007f68fffff3b3;
    assign coff[252 ] = 64'h00007f67fffff3a6;
    assign coff[253 ] = 64'h00007f66fffff39a;
    assign coff[254 ] = 64'h00007f65fffff38d;
    assign coff[255 ] = 64'h00007f63fffff381;
    assign coff[256 ] = 64'h00007f62fffff374;
    assign coff[257 ] = 64'h00007f61fffff368;
    assign coff[258 ] = 64'h00007f60fffff35b;
    assign coff[259 ] = 64'h00007f5efffff34f;
    assign coff[260 ] = 64'h00007f5dfffff342;
    assign coff[261 ] = 64'h00007f5cfffff336;
    assign coff[262 ] = 64'h00007f5bfffff329;
    assign coff[263 ] = 64'h00007f59fffff31d;
    assign coff[264 ] = 64'h00007f58fffff310;
    assign coff[265 ] = 64'h00007f57fffff304;
    assign coff[266 ] = 64'h00007f56fffff2f7;
    assign coff[267 ] = 64'h00007f54fffff2eb;
    assign coff[268 ] = 64'h00007f53fffff2de;
    assign coff[269 ] = 64'h00007f52fffff2d2;
    assign coff[270 ] = 64'h00007f50fffff2c5;
    assign coff[271 ] = 64'h00007f4ffffff2b9;
    assign coff[272 ] = 64'h00007f4efffff2ac;
    assign coff[273 ] = 64'h00007f4dfffff2a0;
    assign coff[274 ] = 64'h00007f4bfffff293;
    assign coff[275 ] = 64'h00007f4afffff287;
    assign coff[276 ] = 64'h00007f49fffff27a;
    assign coff[277 ] = 64'h00007f47fffff26e;
    assign coff[278 ] = 64'h00007f46fffff261;
    assign coff[279 ] = 64'h00007f45fffff255;
    assign coff[280 ] = 64'h00007f43fffff248;
    assign coff[281 ] = 64'h00007f42fffff23c;
    assign coff[282 ] = 64'h00007f41fffff22f;
    assign coff[283 ] = 64'h00007f3ffffff223;
    assign coff[284 ] = 64'h00007f3efffff216;
    assign coff[285 ] = 64'h00007f3cfffff20a;
    assign coff[286 ] = 64'h00007f3bfffff1fd;
    assign coff[287 ] = 64'h00007f3afffff1f1;
    assign coff[288 ] = 64'h00007f38fffff1e4;
    assign coff[289 ] = 64'h00007f37fffff1d8;
    assign coff[290 ] = 64'h00007f36fffff1cb;
    assign coff[291 ] = 64'h00007f34fffff1bf;
    assign coff[292 ] = 64'h00007f33fffff1b2;
    assign coff[293 ] = 64'h00007f31fffff1a6;
    assign coff[294 ] = 64'h00007f30fffff199;
    assign coff[295 ] = 64'h00007f2ffffff18d;
    assign coff[296 ] = 64'h00007f2dfffff180;
    assign coff[297 ] = 64'h00007f2cfffff174;
    assign coff[298 ] = 64'h00007f2afffff167;
    assign coff[299 ] = 64'h00007f29fffff15b;
    assign coff[300 ] = 64'h00007f27fffff14e;
    assign coff[301 ] = 64'h00007f26fffff142;
    assign coff[302 ] = 64'h00007f24fffff135;
    assign coff[303 ] = 64'h00007f23fffff129;
    assign coff[304 ] = 64'h00007f22fffff11c;
    assign coff[305 ] = 64'h00007f20fffff110;
    assign coff[306 ] = 64'h00007f1ffffff104;
    assign coff[307 ] = 64'h00007f1dfffff0f7;
    assign coff[308 ] = 64'h00007f1cfffff0eb;
    assign coff[309 ] = 64'h00007f1afffff0de;
    assign coff[310 ] = 64'h00007f19fffff0d2;
    assign coff[311 ] = 64'h00007f17fffff0c5;
    assign coff[312 ] = 64'h00007f16fffff0b9;
    assign coff[313 ] = 64'h00007f14fffff0ac;
    assign coff[314 ] = 64'h00007f13fffff0a0;
    assign coff[315 ] = 64'h00007f11fffff093;
    assign coff[316 ] = 64'h00007f10fffff087;
    assign coff[317 ] = 64'h00007f0efffff07a;
    assign coff[318 ] = 64'h00007f0dfffff06e;
    assign coff[319 ] = 64'h00007f0bfffff061;
    assign coff[320 ] = 64'h00007f0afffff055;
    assign coff[321 ] = 64'h00007f08fffff048;
    assign coff[322 ] = 64'h00007f06fffff03c;
    assign coff[323 ] = 64'h00007f05fffff02f;
    assign coff[324 ] = 64'h00007f03fffff023;
    assign coff[325 ] = 64'h00007f02fffff016;
    assign coff[326 ] = 64'h00007f00fffff00a;
    assign coff[327 ] = 64'h00007effffffeffe;
    assign coff[328 ] = 64'h00007efdffffeff1;
    assign coff[329 ] = 64'h00007efcffffefe5;
    assign coff[330 ] = 64'h00007efaffffefd8;
    assign coff[331 ] = 64'h00007ef8ffffefcc;
    assign coff[332 ] = 64'h00007ef7ffffefbf;
    assign coff[333 ] = 64'h00007ef5ffffefb3;
    assign coff[334 ] = 64'h00007ef4ffffefa6;
    assign coff[335 ] = 64'h00007ef2ffffef9a;
    assign coff[336 ] = 64'h00007ef0ffffef8d;
    assign coff[337 ] = 64'h00007eefffffef81;
    assign coff[338 ] = 64'h00007eedffffef74;
    assign coff[339 ] = 64'h00007eebffffef68;
    assign coff[340 ] = 64'h00007eeaffffef5c;
    assign coff[341 ] = 64'h00007ee8ffffef4f;
    assign coff[342 ] = 64'h00007ee7ffffef43;
    assign coff[343 ] = 64'h00007ee5ffffef36;
    assign coff[344 ] = 64'h00007ee3ffffef2a;
    assign coff[345 ] = 64'h00007ee2ffffef1d;
    assign coff[346 ] = 64'h00007ee0ffffef11;
    assign coff[347 ] = 64'h00007edeffffef04;
    assign coff[348 ] = 64'h00007eddffffeef8;
    assign coff[349 ] = 64'h00007edbffffeeeb;
    assign coff[350 ] = 64'h00007ed9ffffeedf;
    assign coff[351 ] = 64'h00007ed8ffffeed3;
    assign coff[352 ] = 64'h00007ed6ffffeec6;
    assign coff[353 ] = 64'h00007ed4ffffeeba;
    assign coff[354 ] = 64'h00007ed3ffffeead;
    assign coff[355 ] = 64'h00007ed1ffffeea1;
    assign coff[356 ] = 64'h00007ecfffffee94;
    assign coff[357 ] = 64'h00007ecdffffee88;
    assign coff[358 ] = 64'h00007eccffffee7b;
    assign coff[359 ] = 64'h00007ecaffffee6f;
    assign coff[360 ] = 64'h00007ec8ffffee62;
    assign coff[361 ] = 64'h00007ec6ffffee56;
    assign coff[362 ] = 64'h00007ec5ffffee4a;
    assign coff[363 ] = 64'h00007ec3ffffee3d;
    assign coff[364 ] = 64'h00007ec1ffffee31;
    assign coff[365 ] = 64'h00007ec0ffffee24;
    assign coff[366 ] = 64'h00007ebeffffee18;
    assign coff[367 ] = 64'h00007ebcffffee0b;
    assign coff[368 ] = 64'h00007ebaffffedff;
    assign coff[369 ] = 64'h00007eb8ffffedf2;
    assign coff[370 ] = 64'h00007eb7ffffede6;
    assign coff[371 ] = 64'h00007eb5ffffedda;
    assign coff[372 ] = 64'h00007eb3ffffedcd;
    assign coff[373 ] = 64'h00007eb1ffffedc1;
    assign coff[374 ] = 64'h00007eb0ffffedb4;
    assign coff[375 ] = 64'h00007eaeffffeda8;
    assign coff[376 ] = 64'h00007eacffffed9b;
    assign coff[377 ] = 64'h00007eaaffffed8f;
    assign coff[378 ] = 64'h00007ea8ffffed83;
    assign coff[379 ] = 64'h00007ea6ffffed76;
    assign coff[380 ] = 64'h00007ea5ffffed6a;
    assign coff[381 ] = 64'h00007ea3ffffed5d;
    assign coff[382 ] = 64'h00007ea1ffffed51;
    assign coff[383 ] = 64'h00007e9fffffed44;
    assign coff[384 ] = 64'h00007e9dffffed38;
    assign coff[385 ] = 64'h00007e9bffffed2c;
    assign coff[386 ] = 64'h00007e9affffed1f;
    assign coff[387 ] = 64'h00007e98ffffed13;
    assign coff[388 ] = 64'h00007e96ffffed06;
    assign coff[389 ] = 64'h00007e94ffffecfa;
    assign coff[390 ] = 64'h00007e92ffffeced;
    assign coff[391 ] = 64'h00007e90ffffece1;
    assign coff[392 ] = 64'h00007e8effffecd5;
    assign coff[393 ] = 64'h00007e8dffffecc8;
    assign coff[394 ] = 64'h00007e8bffffecbc;
    assign coff[395 ] = 64'h00007e89ffffecaf;
    assign coff[396 ] = 64'h00007e87ffffeca3;
    assign coff[397 ] = 64'h00007e85ffffec96;
    assign coff[398 ] = 64'h00007e83ffffec8a;
    assign coff[399 ] = 64'h00007e81ffffec7e;
    assign coff[400 ] = 64'h00007e7fffffec71;
    assign coff[401 ] = 64'h00007e7dffffec65;
    assign coff[402 ] = 64'h00007e7bffffec58;
    assign coff[403 ] = 64'h00007e79ffffec4c;
    assign coff[404 ] = 64'h00007e78ffffec3f;
    assign coff[405 ] = 64'h00007e76ffffec33;
    assign coff[406 ] = 64'h00007e74ffffec27;
    assign coff[407 ] = 64'h00007e72ffffec1a;
    assign coff[408 ] = 64'h00007e70ffffec0e;
    assign coff[409 ] = 64'h00007e6effffec01;
    assign coff[410 ] = 64'h00007e6cffffebf5;
    assign coff[411 ] = 64'h00007e6affffebe9;
    assign coff[412 ] = 64'h00007e68ffffebdc;
    assign coff[413 ] = 64'h00007e66ffffebd0;
    assign coff[414 ] = 64'h00007e64ffffebc3;
    assign coff[415 ] = 64'h00007e62ffffebb7;
    assign coff[416 ] = 64'h00007e60ffffebab;
    assign coff[417 ] = 64'h00007e5effffeb9e;
    assign coff[418 ] = 64'h00007e5cffffeb92;
    assign coff[419 ] = 64'h00007e5affffeb85;
    assign coff[420 ] = 64'h00007e58ffffeb79;
    assign coff[421 ] = 64'h00007e56ffffeb6d;
    assign coff[422 ] = 64'h00007e54ffffeb60;
    assign coff[423 ] = 64'h00007e52ffffeb54;
    assign coff[424 ] = 64'h00007e50ffffeb47;
    assign coff[425 ] = 64'h00007e4effffeb3b;
    assign coff[426 ] = 64'h00007e4cffffeb2f;
    assign coff[427 ] = 64'h00007e4affffeb22;
    assign coff[428 ] = 64'h00007e48ffffeb16;
    assign coff[429 ] = 64'h00007e46ffffeb09;
    assign coff[430 ] = 64'h00007e43ffffeafd;
    assign coff[431 ] = 64'h00007e41ffffeaf1;
    assign coff[432 ] = 64'h00007e3fffffeae4;
    assign coff[433 ] = 64'h00007e3dffffead8;
    assign coff[434 ] = 64'h00007e3bffffeacb;
    assign coff[435 ] = 64'h00007e39ffffeabf;
    assign coff[436 ] = 64'h00007e37ffffeab3;
    assign coff[437 ] = 64'h00007e35ffffeaa6;
    assign coff[438 ] = 64'h00007e33ffffea9a;
    assign coff[439 ] = 64'h00007e31ffffea8d;
    assign coff[440 ] = 64'h00007e2fffffea81;
    assign coff[441 ] = 64'h00007e2dffffea75;
    assign coff[442 ] = 64'h00007e2affffea68;
    assign coff[443 ] = 64'h00007e28ffffea5c;
    assign coff[444 ] = 64'h00007e26ffffea4f;
    assign coff[445 ] = 64'h00007e24ffffea43;
    assign coff[446 ] = 64'h00007e22ffffea37;
    assign coff[447 ] = 64'h00007e20ffffea2a;
    assign coff[448 ] = 64'h00007e1effffea1e;
    assign coff[449 ] = 64'h00007e1bffffea12;
    assign coff[450 ] = 64'h00007e19ffffea05;
    assign coff[451 ] = 64'h00007e17ffffe9f9;
    assign coff[452 ] = 64'h00007e15ffffe9ec;
    assign coff[453 ] = 64'h00007e13ffffe9e0;
    assign coff[454 ] = 64'h00007e11ffffe9d4;
    assign coff[455 ] = 64'h00007e0effffe9c7;
    assign coff[456 ] = 64'h00007e0cffffe9bb;
    assign coff[457 ] = 64'h00007e0affffe9af;
    assign coff[458 ] = 64'h00007e08ffffe9a2;
    assign coff[459 ] = 64'h00007e06ffffe996;
    assign coff[460 ] = 64'h00007e03ffffe989;
    assign coff[461 ] = 64'h00007e01ffffe97d;
    assign coff[462 ] = 64'h00007dffffffe971;
    assign coff[463 ] = 64'h00007dfdffffe964;
    assign coff[464 ] = 64'h00007dfbffffe958;
    assign coff[465 ] = 64'h00007df8ffffe94c;
    assign coff[466 ] = 64'h00007df6ffffe93f;
    assign coff[467 ] = 64'h00007df4ffffe933;
    assign coff[468 ] = 64'h00007df2ffffe926;
    assign coff[469 ] = 64'h00007defffffe91a;
    assign coff[470 ] = 64'h00007dedffffe90e;
    assign coff[471 ] = 64'h00007debffffe901;
    assign coff[472 ] = 64'h00007de9ffffe8f5;
    assign coff[473 ] = 64'h00007de6ffffe8e9;
    assign coff[474 ] = 64'h00007de4ffffe8dc;
    assign coff[475 ] = 64'h00007de2ffffe8d0;
    assign coff[476 ] = 64'h00007de0ffffe8c4;
    assign coff[477 ] = 64'h00007dddffffe8b7;
    assign coff[478 ] = 64'h00007ddbffffe8ab;
    assign coff[479 ] = 64'h00007dd9ffffe89f;
    assign coff[480 ] = 64'h00007dd6ffffe892;
    assign coff[481 ] = 64'h00007dd4ffffe886;
    assign coff[482 ] = 64'h00007dd2ffffe879;
    assign coff[483 ] = 64'h00007dcfffffe86d;
    assign coff[484 ] = 64'h00007dcdffffe861;
    assign coff[485 ] = 64'h00007dcbffffe854;
    assign coff[486 ] = 64'h00007dc9ffffe848;
    assign coff[487 ] = 64'h00007dc6ffffe83c;
    assign coff[488 ] = 64'h00007dc4ffffe82f;
    assign coff[489 ] = 64'h00007dc2ffffe823;
    assign coff[490 ] = 64'h00007dbfffffe817;
    assign coff[491 ] = 64'h00007dbdffffe80a;
    assign coff[492 ] = 64'h00007dbaffffe7fe;
    assign coff[493 ] = 64'h00007db8ffffe7f2;
    assign coff[494 ] = 64'h00007db6ffffe7e5;
    assign coff[495 ] = 64'h00007db3ffffe7d9;
    assign coff[496 ] = 64'h00007db1ffffe7cd;
    assign coff[497 ] = 64'h00007dafffffe7c0;
    assign coff[498 ] = 64'h00007dacffffe7b4;
    assign coff[499 ] = 64'h00007daaffffe7a8;
    assign coff[500 ] = 64'h00007da7ffffe79b;
    assign coff[501 ] = 64'h00007da5ffffe78f;
    assign coff[502 ] = 64'h00007da3ffffe783;
    assign coff[503 ] = 64'h00007da0ffffe776;
    assign coff[504 ] = 64'h00007d9effffe76a;
    assign coff[505 ] = 64'h00007d9bffffe75e;
    assign coff[506 ] = 64'h00007d99ffffe751;
    assign coff[507 ] = 64'h00007d97ffffe745;
    assign coff[508 ] = 64'h00007d94ffffe739;
    assign coff[509 ] = 64'h00007d92ffffe72c;
    assign coff[510 ] = 64'h00007d8fffffe720;
    assign coff[511 ] = 64'h00007d8dffffe714;
    assign coff[512 ] = 64'h00007d8affffe707;
    assign coff[513 ] = 64'h00007d88ffffe6fb;
    assign coff[514 ] = 64'h00007d85ffffe6ef;
    assign coff[515 ] = 64'h00007d83ffffe6e2;
    assign coff[516 ] = 64'h00007d81ffffe6d6;
    assign coff[517 ] = 64'h00007d7effffe6ca;
    assign coff[518 ] = 64'h00007d7cffffe6bd;
    assign coff[519 ] = 64'h00007d79ffffe6b1;
    assign coff[520 ] = 64'h00007d77ffffe6a5;
    assign coff[521 ] = 64'h00007d74ffffe698;
    assign coff[522 ] = 64'h00007d72ffffe68c;
    assign coff[523 ] = 64'h00007d6fffffe680;
    assign coff[524 ] = 64'h00007d6dffffe673;
    assign coff[525 ] = 64'h00007d6affffe667;
    assign coff[526 ] = 64'h00007d68ffffe65b;
    assign coff[527 ] = 64'h00007d65ffffe64f;
    assign coff[528 ] = 64'h00007d63ffffe642;
    assign coff[529 ] = 64'h00007d60ffffe636;
    assign coff[530 ] = 64'h00007d5dffffe62a;
    assign coff[531 ] = 64'h00007d5bffffe61d;
    assign coff[532 ] = 64'h00007d58ffffe611;
    assign coff[533 ] = 64'h00007d56ffffe605;
    assign coff[534 ] = 64'h00007d53ffffe5f8;
    assign coff[535 ] = 64'h00007d51ffffe5ec;
    assign coff[536 ] = 64'h00007d4effffe5e0;
    assign coff[537 ] = 64'h00007d4cffffe5d3;
    assign coff[538 ] = 64'h00007d49ffffe5c7;
    assign coff[539 ] = 64'h00007d46ffffe5bb;
    assign coff[540 ] = 64'h00007d44ffffe5af;
    assign coff[541 ] = 64'h00007d41ffffe5a2;
    assign coff[542 ] = 64'h00007d3fffffe596;
    assign coff[543 ] = 64'h00007d3cffffe58a;
    assign coff[544 ] = 64'h00007d3affffe57d;
    assign coff[545 ] = 64'h00007d37ffffe571;
    assign coff[546 ] = 64'h00007d34ffffe565;
    assign coff[547 ] = 64'h00007d32ffffe558;
    assign coff[548 ] = 64'h00007d2fffffe54c;
    assign coff[549 ] = 64'h00007d2cffffe540;
    assign coff[550 ] = 64'h00007d2affffe534;
    assign coff[551 ] = 64'h00007d27ffffe527;
    assign coff[552 ] = 64'h00007d25ffffe51b;
    assign coff[553 ] = 64'h00007d22ffffe50f;
    assign coff[554 ] = 64'h00007d1fffffe502;
    assign coff[555 ] = 64'h00007d1dffffe4f6;
    assign coff[556 ] = 64'h00007d1affffe4ea;
    assign coff[557 ] = 64'h00007d17ffffe4de;
    assign coff[558 ] = 64'h00007d15ffffe4d1;
    assign coff[559 ] = 64'h00007d12ffffe4c5;
    assign coff[560 ] = 64'h00007d0fffffe4b9;
    assign coff[561 ] = 64'h00007d0dffffe4ad;
    assign coff[562 ] = 64'h00007d0affffe4a0;
    assign coff[563 ] = 64'h00007d07ffffe494;
    assign coff[564 ] = 64'h00007d05ffffe488;
    assign coff[565 ] = 64'h00007d02ffffe47b;
    assign coff[566 ] = 64'h00007cffffffe46f;
    assign coff[567 ] = 64'h00007cfcffffe463;
    assign coff[568 ] = 64'h00007cfaffffe457;
    assign coff[569 ] = 64'h00007cf7ffffe44a;
    assign coff[570 ] = 64'h00007cf4ffffe43e;
    assign coff[571 ] = 64'h00007cf2ffffe432;
    assign coff[572 ] = 64'h00007cefffffe426;
    assign coff[573 ] = 64'h00007cecffffe419;
    assign coff[574 ] = 64'h00007ce9ffffe40d;
    assign coff[575 ] = 64'h00007ce7ffffe401;
    assign coff[576 ] = 64'h00007ce4ffffe3f4;
    assign coff[577 ] = 64'h00007ce1ffffe3e8;
    assign coff[578 ] = 64'h00007cdeffffe3dc;
    assign coff[579 ] = 64'h00007cdcffffe3d0;
    assign coff[580 ] = 64'h00007cd9ffffe3c3;
    assign coff[581 ] = 64'h00007cd6ffffe3b7;
    assign coff[582 ] = 64'h00007cd3ffffe3ab;
    assign coff[583 ] = 64'h00007cd0ffffe39f;
    assign coff[584 ] = 64'h00007cceffffe392;
    assign coff[585 ] = 64'h00007ccbffffe386;
    assign coff[586 ] = 64'h00007cc8ffffe37a;
    assign coff[587 ] = 64'h00007cc5ffffe36e;
    assign coff[588 ] = 64'h00007cc2ffffe361;
    assign coff[589 ] = 64'h00007cc0ffffe355;
    assign coff[590 ] = 64'h00007cbdffffe349;
    assign coff[591 ] = 64'h00007cbaffffe33d;
    assign coff[592 ] = 64'h00007cb7ffffe330;
    assign coff[593 ] = 64'h00007cb4ffffe324;
    assign coff[594 ] = 64'h00007cb1ffffe318;
    assign coff[595 ] = 64'h00007cafffffe30c;
    assign coff[596 ] = 64'h00007cacffffe2ff;
    assign coff[597 ] = 64'h00007ca9ffffe2f3;
    assign coff[598 ] = 64'h00007ca6ffffe2e7;
    assign coff[599 ] = 64'h00007ca3ffffe2db;
    assign coff[600 ] = 64'h00007ca0ffffe2cf;
    assign coff[601 ] = 64'h00007c9effffe2c2;
    assign coff[602 ] = 64'h00007c9bffffe2b6;
    assign coff[603 ] = 64'h00007c98ffffe2aa;
    assign coff[604 ] = 64'h00007c95ffffe29e;
    assign coff[605 ] = 64'h00007c92ffffe291;
    assign coff[606 ] = 64'h00007c8fffffe285;
    assign coff[607 ] = 64'h00007c8cffffe279;
    assign coff[608 ] = 64'h00007c89ffffe26d;
    assign coff[609 ] = 64'h00007c86ffffe260;
    assign coff[610 ] = 64'h00007c83ffffe254;
    assign coff[611 ] = 64'h00007c81ffffe248;
    assign coff[612 ] = 64'h00007c7effffe23c;
    assign coff[613 ] = 64'h00007c7bffffe230;
    assign coff[614 ] = 64'h00007c78ffffe223;
    assign coff[615 ] = 64'h00007c75ffffe217;
    assign coff[616 ] = 64'h00007c72ffffe20b;
    assign coff[617 ] = 64'h00007c6fffffe1ff;
    assign coff[618 ] = 64'h00007c6cffffe1f2;
    assign coff[619 ] = 64'h00007c69ffffe1e6;
    assign coff[620 ] = 64'h00007c66ffffe1da;
    assign coff[621 ] = 64'h00007c63ffffe1ce;
    assign coff[622 ] = 64'h00007c60ffffe1c2;
    assign coff[623 ] = 64'h00007c5dffffe1b5;
    assign coff[624 ] = 64'h00007c5affffe1a9;
    assign coff[625 ] = 64'h00007c57ffffe19d;
    assign coff[626 ] = 64'h00007c54ffffe191;
    assign coff[627 ] = 64'h00007c51ffffe185;
    assign coff[628 ] = 64'h00007c4effffe178;
    assign coff[629 ] = 64'h00007c4bffffe16c;
    assign coff[630 ] = 64'h00007c48ffffe160;
    assign coff[631 ] = 64'h00007c45ffffe154;
    assign coff[632 ] = 64'h00007c42ffffe148;
    assign coff[633 ] = 64'h00007c3fffffe13b;
    assign coff[634 ] = 64'h00007c3cffffe12f;
    assign coff[635 ] = 64'h00007c39ffffe123;
    assign coff[636 ] = 64'h00007c36ffffe117;
    assign coff[637 ] = 64'h00007c33ffffe10b;
    assign coff[638 ] = 64'h00007c30ffffe0fe;
    assign coff[639 ] = 64'h00007c2dffffe0f2;
    assign coff[640 ] = 64'h00007c2affffe0e6;
    assign coff[641 ] = 64'h00007c27ffffe0da;
    assign coff[642 ] = 64'h00007c24ffffe0ce;
    assign coff[643 ] = 64'h00007c21ffffe0c1;
    assign coff[644 ] = 64'h00007c1effffe0b5;
    assign coff[645 ] = 64'h00007c1bffffe0a9;
    assign coff[646 ] = 64'h00007c18ffffe09d;
    assign coff[647 ] = 64'h00007c14ffffe091;
    assign coff[648 ] = 64'h00007c11ffffe085;
    assign coff[649 ] = 64'h00007c0effffe078;
    assign coff[650 ] = 64'h00007c0bffffe06c;
    assign coff[651 ] = 64'h00007c08ffffe060;
    assign coff[652 ] = 64'h00007c05ffffe054;
    assign coff[653 ] = 64'h00007c02ffffe048;
    assign coff[654 ] = 64'h00007bffffffe03b;
    assign coff[655 ] = 64'h00007bfcffffe02f;
    assign coff[656 ] = 64'h00007bf9ffffe023;
    assign coff[657 ] = 64'h00007bf5ffffe017;
    assign coff[658 ] = 64'h00007bf2ffffe00b;
    assign coff[659 ] = 64'h00007befffffdfff;
    assign coff[660 ] = 64'h00007becffffdff2;
    assign coff[661 ] = 64'h00007be9ffffdfe6;
    assign coff[662 ] = 64'h00007be6ffffdfda;
    assign coff[663 ] = 64'h00007be3ffffdfce;
    assign coff[664 ] = 64'h00007bdfffffdfc2;
    assign coff[665 ] = 64'h00007bdcffffdfb6;
    assign coff[666 ] = 64'h00007bd9ffffdfa9;
    assign coff[667 ] = 64'h00007bd6ffffdf9d;
    assign coff[668 ] = 64'h00007bd3ffffdf91;
    assign coff[669 ] = 64'h00007bcfffffdf85;
    assign coff[670 ] = 64'h00007bccffffdf79;
    assign coff[671 ] = 64'h00007bc9ffffdf6d;
    assign coff[672 ] = 64'h00007bc6ffffdf61;
    assign coff[673 ] = 64'h00007bc3ffffdf54;
    assign coff[674 ] = 64'h00007bbfffffdf48;
    assign coff[675 ] = 64'h00007bbcffffdf3c;
    assign coff[676 ] = 64'h00007bb9ffffdf30;
    assign coff[677 ] = 64'h00007bb6ffffdf24;
    assign coff[678 ] = 64'h00007bb3ffffdf18;
    assign coff[679 ] = 64'h00007bafffffdf0c;
    assign coff[680 ] = 64'h00007bacffffdeff;
    assign coff[681 ] = 64'h00007ba9ffffdef3;
    assign coff[682 ] = 64'h00007ba6ffffdee7;
    assign coff[683 ] = 64'h00007ba2ffffdedb;
    assign coff[684 ] = 64'h00007b9fffffdecf;
    assign coff[685 ] = 64'h00007b9cffffdec3;
    assign coff[686 ] = 64'h00007b99ffffdeb7;
    assign coff[687 ] = 64'h00007b95ffffdeaa;
    assign coff[688 ] = 64'h00007b92ffffde9e;
    assign coff[689 ] = 64'h00007b8fffffde92;
    assign coff[690 ] = 64'h00007b8bffffde86;
    assign coff[691 ] = 64'h00007b88ffffde7a;
    assign coff[692 ] = 64'h00007b85ffffde6e;
    assign coff[693 ] = 64'h00007b82ffffde62;
    assign coff[694 ] = 64'h00007b7effffde56;
    assign coff[695 ] = 64'h00007b7bffffde49;
    assign coff[696 ] = 64'h00007b78ffffde3d;
    assign coff[697 ] = 64'h00007b74ffffde31;
    assign coff[698 ] = 64'h00007b71ffffde25;
    assign coff[699 ] = 64'h00007b6effffde19;
    assign coff[700 ] = 64'h00007b6affffde0d;
    assign coff[701 ] = 64'h00007b67ffffde01;
    assign coff[702 ] = 64'h00007b64ffffddf5;
    assign coff[703 ] = 64'h00007b60ffffdde8;
    assign coff[704 ] = 64'h00007b5dffffdddc;
    assign coff[705 ] = 64'h00007b5affffddd0;
    assign coff[706 ] = 64'h00007b56ffffddc4;
    assign coff[707 ] = 64'h00007b53ffffddb8;
    assign coff[708 ] = 64'h00007b50ffffddac;
    assign coff[709 ] = 64'h00007b4cffffdda0;
    assign coff[710 ] = 64'h00007b49ffffdd94;
    assign coff[711 ] = 64'h00007b45ffffdd88;
    assign coff[712 ] = 64'h00007b42ffffdd7c;
    assign coff[713 ] = 64'h00007b3fffffdd6f;
    assign coff[714 ] = 64'h00007b3bffffdd63;
    assign coff[715 ] = 64'h00007b38ffffdd57;
    assign coff[716 ] = 64'h00007b34ffffdd4b;
    assign coff[717 ] = 64'h00007b31ffffdd3f;
    assign coff[718 ] = 64'h00007b2effffdd33;
    assign coff[719 ] = 64'h00007b2affffdd27;
    assign coff[720 ] = 64'h00007b27ffffdd1b;
    assign coff[721 ] = 64'h00007b23ffffdd0f;
    assign coff[722 ] = 64'h00007b20ffffdd03;
    assign coff[723 ] = 64'h00007b1cffffdcf6;
    assign coff[724 ] = 64'h00007b19ffffdcea;
    assign coff[725 ] = 64'h00007b16ffffdcde;
    assign coff[726 ] = 64'h00007b12ffffdcd2;
    assign coff[727 ] = 64'h00007b0fffffdcc6;
    assign coff[728 ] = 64'h00007b0bffffdcba;
    assign coff[729 ] = 64'h00007b08ffffdcae;
    assign coff[730 ] = 64'h00007b04ffffdca2;
    assign coff[731 ] = 64'h00007b01ffffdc96;
    assign coff[732 ] = 64'h00007afdffffdc8a;
    assign coff[733 ] = 64'h00007afaffffdc7e;
    assign coff[734 ] = 64'h00007af6ffffdc72;
    assign coff[735 ] = 64'h00007af3ffffdc66;
    assign coff[736 ] = 64'h00007aefffffdc59;
    assign coff[737 ] = 64'h00007aecffffdc4d;
    assign coff[738 ] = 64'h00007ae8ffffdc41;
    assign coff[739 ] = 64'h00007ae5ffffdc35;
    assign coff[740 ] = 64'h00007ae1ffffdc29;
    assign coff[741 ] = 64'h00007adeffffdc1d;
    assign coff[742 ] = 64'h00007adaffffdc11;
    assign coff[743 ] = 64'h00007ad7ffffdc05;
    assign coff[744 ] = 64'h00007ad3ffffdbf9;
    assign coff[745 ] = 64'h00007ad0ffffdbed;
    assign coff[746 ] = 64'h00007accffffdbe1;
    assign coff[747 ] = 64'h00007ac9ffffdbd5;
    assign coff[748 ] = 64'h00007ac5ffffdbc9;
    assign coff[749 ] = 64'h00007ac1ffffdbbd;
    assign coff[750 ] = 64'h00007abeffffdbb1;
    assign coff[751 ] = 64'h00007abaffffdba5;
    assign coff[752 ] = 64'h00007ab7ffffdb99;
    assign coff[753 ] = 64'h00007ab3ffffdb8c;
    assign coff[754 ] = 64'h00007ab0ffffdb80;
    assign coff[755 ] = 64'h00007aacffffdb74;
    assign coff[756 ] = 64'h00007aa8ffffdb68;
    assign coff[757 ] = 64'h00007aa5ffffdb5c;
    assign coff[758 ] = 64'h00007aa1ffffdb50;
    assign coff[759 ] = 64'h00007a9effffdb44;
    assign coff[760 ] = 64'h00007a9affffdb38;
    assign coff[761 ] = 64'h00007a96ffffdb2c;
    assign coff[762 ] = 64'h00007a93ffffdb20;
    assign coff[763 ] = 64'h00007a8fffffdb14;
    assign coff[764 ] = 64'h00007a8cffffdb08;
    assign coff[765 ] = 64'h00007a88ffffdafc;
    assign coff[766 ] = 64'h00007a84ffffdaf0;
    assign coff[767 ] = 64'h00007a81ffffdae4;
    assign coff[768 ] = 64'h00007a7dffffdad8;
    assign coff[769 ] = 64'h00007a79ffffdacc;
    assign coff[770 ] = 64'h00007a76ffffdac0;
    assign coff[771 ] = 64'h00007a72ffffdab4;
    assign coff[772 ] = 64'h00007a6effffdaa8;
    assign coff[773 ] = 64'h00007a6bffffda9c;
    assign coff[774 ] = 64'h00007a67ffffda90;
    assign coff[775 ] = 64'h00007a63ffffda84;
    assign coff[776 ] = 64'h00007a60ffffda78;
    assign coff[777 ] = 64'h00007a5cffffda6c;
    assign coff[778 ] = 64'h00007a58ffffda60;
    assign coff[779 ] = 64'h00007a55ffffda54;
    assign coff[780 ] = 64'h00007a51ffffda48;
    assign coff[781 ] = 64'h00007a4dffffda3c;
    assign coff[782 ] = 64'h00007a49ffffda30;
    assign coff[783 ] = 64'h00007a46ffffda24;
    assign coff[784 ] = 64'h00007a42ffffda18;
    assign coff[785 ] = 64'h00007a3effffda0c;
    assign coff[786 ] = 64'h00007a3bffffda00;
    assign coff[787 ] = 64'h00007a37ffffd9f4;
    assign coff[788 ] = 64'h00007a33ffffd9e8;
    assign coff[789 ] = 64'h00007a2fffffd9dc;
    assign coff[790 ] = 64'h00007a2cffffd9d0;
    assign coff[791 ] = 64'h00007a28ffffd9c4;
    assign coff[792 ] = 64'h00007a24ffffd9b8;
    assign coff[793 ] = 64'h00007a20ffffd9ac;
    assign coff[794 ] = 64'h00007a1dffffd9a0;
    assign coff[795 ] = 64'h00007a19ffffd994;
    assign coff[796 ] = 64'h00007a15ffffd988;
    assign coff[797 ] = 64'h00007a11ffffd97c;
    assign coff[798 ] = 64'h00007a0effffd970;
    assign coff[799 ] = 64'h00007a0affffd964;
    assign coff[800 ] = 64'h00007a06ffffd958;
    assign coff[801 ] = 64'h00007a02ffffd94c;
    assign coff[802 ] = 64'h000079feffffd940;
    assign coff[803 ] = 64'h000079fbffffd934;
    assign coff[804 ] = 64'h000079f7ffffd928;
    assign coff[805 ] = 64'h000079f3ffffd91c;
    assign coff[806 ] = 64'h000079efffffd910;
    assign coff[807 ] = 64'h000079ebffffd904;
    assign coff[808 ] = 64'h000079e7ffffd8f8;
    assign coff[809 ] = 64'h000079e4ffffd8ec;
    assign coff[810 ] = 64'h000079e0ffffd8e0;
    assign coff[811 ] = 64'h000079dcffffd8d4;
    assign coff[812 ] = 64'h000079d8ffffd8c8;
    assign coff[813 ] = 64'h000079d4ffffd8bc;
    assign coff[814 ] = 64'h000079d0ffffd8b0;
    assign coff[815 ] = 64'h000079ccffffd8a4;
    assign coff[816 ] = 64'h000079c9ffffd898;
    assign coff[817 ] = 64'h000079c5ffffd88c;
    assign coff[818 ] = 64'h000079c1ffffd880;
    assign coff[819 ] = 64'h000079bdffffd875;
    assign coff[820 ] = 64'h000079b9ffffd869;
    assign coff[821 ] = 64'h000079b5ffffd85d;
    assign coff[822 ] = 64'h000079b1ffffd851;
    assign coff[823 ] = 64'h000079adffffd845;
    assign coff[824 ] = 64'h000079aaffffd839;
    assign coff[825 ] = 64'h000079a6ffffd82d;
    assign coff[826 ] = 64'h000079a2ffffd821;
    assign coff[827 ] = 64'h0000799effffd815;
    assign coff[828 ] = 64'h0000799affffd809;
    assign coff[829 ] = 64'h00007996ffffd7fd;
    assign coff[830 ] = 64'h00007992ffffd7f1;
    assign coff[831 ] = 64'h0000798effffd7e5;
    assign coff[832 ] = 64'h0000798affffd7d9;
    assign coff[833 ] = 64'h00007986ffffd7cd;
    assign coff[834 ] = 64'h00007982ffffd7c1;
    assign coff[835 ] = 64'h0000797effffd7b5;
    assign coff[836 ] = 64'h0000797affffd7aa;
    assign coff[837 ] = 64'h00007976ffffd79e;
    assign coff[838 ] = 64'h00007972ffffd792;
    assign coff[839 ] = 64'h0000796effffd786;
    assign coff[840 ] = 64'h0000796affffd77a;
    assign coff[841 ] = 64'h00007966ffffd76e;
    assign coff[842 ] = 64'h00007962ffffd762;
    assign coff[843 ] = 64'h0000795fffffd756;
    assign coff[844 ] = 64'h0000795bffffd74a;
    assign coff[845 ] = 64'h00007957ffffd73e;
    assign coff[846 ] = 64'h00007953ffffd732;
    assign coff[847 ] = 64'h0000794effffd726;
    assign coff[848 ] = 64'h0000794affffd71b;
    assign coff[849 ] = 64'h00007946ffffd70f;
    assign coff[850 ] = 64'h00007942ffffd703;
    assign coff[851 ] = 64'h0000793effffd6f7;
    assign coff[852 ] = 64'h0000793affffd6eb;
    assign coff[853 ] = 64'h00007936ffffd6df;
    assign coff[854 ] = 64'h00007932ffffd6d3;
    assign coff[855 ] = 64'h0000792effffd6c7;
    assign coff[856 ] = 64'h0000792affffd6bb;
    assign coff[857 ] = 64'h00007926ffffd6af;
    assign coff[858 ] = 64'h00007922ffffd6a4;
    assign coff[859 ] = 64'h0000791effffd698;
    assign coff[860 ] = 64'h0000791affffd68c;
    assign coff[861 ] = 64'h00007916ffffd680;
    assign coff[862 ] = 64'h00007912ffffd674;
    assign coff[863 ] = 64'h0000790effffd668;
    assign coff[864 ] = 64'h0000790affffd65c;
    assign coff[865 ] = 64'h00007906ffffd650;
    assign coff[866 ] = 64'h00007901ffffd644;
    assign coff[867 ] = 64'h000078fdffffd639;
    assign coff[868 ] = 64'h000078f9ffffd62d;
    assign coff[869 ] = 64'h000078f5ffffd621;
    assign coff[870 ] = 64'h000078f1ffffd615;
    assign coff[871 ] = 64'h000078edffffd609;
    assign coff[872 ] = 64'h000078e9ffffd5fd;
    assign coff[873 ] = 64'h000078e5ffffd5f1;
    assign coff[874 ] = 64'h000078e1ffffd5e5;
    assign coff[875 ] = 64'h000078dcffffd5da;
    assign coff[876 ] = 64'h000078d8ffffd5ce;
    assign coff[877 ] = 64'h000078d4ffffd5c2;
    assign coff[878 ] = 64'h000078d0ffffd5b6;
    assign coff[879 ] = 64'h000078ccffffd5aa;
    assign coff[880 ] = 64'h000078c8ffffd59e;
    assign coff[881 ] = 64'h000078c4ffffd592;
    assign coff[882 ] = 64'h000078bfffffd587;
    assign coff[883 ] = 64'h000078bbffffd57b;
    assign coff[884 ] = 64'h000078b7ffffd56f;
    assign coff[885 ] = 64'h000078b3ffffd563;
    assign coff[886 ] = 64'h000078afffffd557;
    assign coff[887 ] = 64'h000078aaffffd54b;
    assign coff[888 ] = 64'h000078a6ffffd53f;
    assign coff[889 ] = 64'h000078a2ffffd534;
    assign coff[890 ] = 64'h0000789effffd528;
    assign coff[891 ] = 64'h0000789affffd51c;
    assign coff[892 ] = 64'h00007895ffffd510;
    assign coff[893 ] = 64'h00007891ffffd504;
    assign coff[894 ] = 64'h0000788dffffd4f8;
    assign coff[895 ] = 64'h00007889ffffd4ed;
    assign coff[896 ] = 64'h00007885ffffd4e1;
    assign coff[897 ] = 64'h00007880ffffd4d5;
    assign coff[898 ] = 64'h0000787cffffd4c9;
    assign coff[899 ] = 64'h00007878ffffd4bd;
    assign coff[900 ] = 64'h00007874ffffd4b1;
    assign coff[901 ] = 64'h0000786fffffd4a6;
    assign coff[902 ] = 64'h0000786bffffd49a;
    assign coff[903 ] = 64'h00007867ffffd48e;
    assign coff[904 ] = 64'h00007863ffffd482;
    assign coff[905 ] = 64'h0000785effffd476;
    assign coff[906 ] = 64'h0000785affffd46b;
    assign coff[907 ] = 64'h00007856ffffd45f;
    assign coff[908 ] = 64'h00007851ffffd453;
    assign coff[909 ] = 64'h0000784dffffd447;
    assign coff[910 ] = 64'h00007849ffffd43b;
    assign coff[911 ] = 64'h00007845ffffd430;
    assign coff[912 ] = 64'h00007840ffffd424;
    assign coff[913 ] = 64'h0000783cffffd418;
    assign coff[914 ] = 64'h00007838ffffd40c;
    assign coff[915 ] = 64'h00007833ffffd400;
    assign coff[916 ] = 64'h0000782fffffd3f4;
    assign coff[917 ] = 64'h0000782bffffd3e9;
    assign coff[918 ] = 64'h00007826ffffd3dd;
    assign coff[919 ] = 64'h00007822ffffd3d1;
    assign coff[920 ] = 64'h0000781effffd3c5;
    assign coff[921 ] = 64'h00007819ffffd3ba;
    assign coff[922 ] = 64'h00007815ffffd3ae;
    assign coff[923 ] = 64'h00007811ffffd3a2;
    assign coff[924 ] = 64'h0000780cffffd396;
    assign coff[925 ] = 64'h00007808ffffd38a;
    assign coff[926 ] = 64'h00007803ffffd37f;
    assign coff[927 ] = 64'h000077ffffffd373;
    assign coff[928 ] = 64'h000077fbffffd367;
    assign coff[929 ] = 64'h000077f6ffffd35b;
    assign coff[930 ] = 64'h000077f2ffffd34f;
    assign coff[931 ] = 64'h000077eeffffd344;
    assign coff[932 ] = 64'h000077e9ffffd338;
    assign coff[933 ] = 64'h000077e5ffffd32c;
    assign coff[934 ] = 64'h000077e0ffffd320;
    assign coff[935 ] = 64'h000077dcffffd315;
    assign coff[936 ] = 64'h000077d8ffffd309;
    assign coff[937 ] = 64'h000077d3ffffd2fd;
    assign coff[938 ] = 64'h000077cfffffd2f1;
    assign coff[939 ] = 64'h000077caffffd2e6;
    assign coff[940 ] = 64'h000077c6ffffd2da;
    assign coff[941 ] = 64'h000077c1ffffd2ce;
    assign coff[942 ] = 64'h000077bdffffd2c2;
    assign coff[943 ] = 64'h000077b9ffffd2b7;
    assign coff[944 ] = 64'h000077b4ffffd2ab;
    assign coff[945 ] = 64'h000077b0ffffd29f;
    assign coff[946 ] = 64'h000077abffffd293;
    assign coff[947 ] = 64'h000077a7ffffd288;
    assign coff[948 ] = 64'h000077a2ffffd27c;
    assign coff[949 ] = 64'h0000779effffd270;
    assign coff[950 ] = 64'h00007799ffffd264;
    assign coff[951 ] = 64'h00007795ffffd259;
    assign coff[952 ] = 64'h00007790ffffd24d;
    assign coff[953 ] = 64'h0000778cffffd241;
    assign coff[954 ] = 64'h00007787ffffd235;
    assign coff[955 ] = 64'h00007783ffffd22a;
    assign coff[956 ] = 64'h0000777effffd21e;
    assign coff[957 ] = 64'h0000777affffd212;
    assign coff[958 ] = 64'h00007775ffffd206;
    assign coff[959 ] = 64'h00007771ffffd1fb;
    assign coff[960 ] = 64'h0000776cffffd1ef;
    assign coff[961 ] = 64'h00007768ffffd1e3;
    assign coff[962 ] = 64'h00007763ffffd1d8;
    assign coff[963 ] = 64'h0000775fffffd1cc;
    assign coff[964 ] = 64'h0000775affffd1c0;
    assign coff[965 ] = 64'h00007756ffffd1b4;
    assign coff[966 ] = 64'h00007751ffffd1a9;
    assign coff[967 ] = 64'h0000774dffffd19d;
    assign coff[968 ] = 64'h00007748ffffd191;
    assign coff[969 ] = 64'h00007743ffffd186;
    assign coff[970 ] = 64'h0000773fffffd17a;
    assign coff[971 ] = 64'h0000773affffd16e;
    assign coff[972 ] = 64'h00007736ffffd162;
    assign coff[973 ] = 64'h00007731ffffd157;
    assign coff[974 ] = 64'h0000772dffffd14b;
    assign coff[975 ] = 64'h00007728ffffd13f;
    assign coff[976 ] = 64'h00007723ffffd134;
    assign coff[977 ] = 64'h0000771fffffd128;
    assign coff[978 ] = 64'h0000771affffd11c;
    assign coff[979 ] = 64'h00007716ffffd111;
    assign coff[980 ] = 64'h00007711ffffd105;
    assign coff[981 ] = 64'h0000770cffffd0f9;
    assign coff[982 ] = 64'h00007708ffffd0ed;
    assign coff[983 ] = 64'h00007703ffffd0e2;
    assign coff[984 ] = 64'h000076feffffd0d6;
    assign coff[985 ] = 64'h000076faffffd0ca;
    assign coff[986 ] = 64'h000076f5ffffd0bf;
    assign coff[987 ] = 64'h000076f1ffffd0b3;
    assign coff[988 ] = 64'h000076ecffffd0a7;
    assign coff[989 ] = 64'h000076e7ffffd09c;
    assign coff[990 ] = 64'h000076e3ffffd090;
    assign coff[991 ] = 64'h000076deffffd084;
    assign coff[992 ] = 64'h000076d9ffffd079;
    assign coff[993 ] = 64'h000076d5ffffd06d;
    assign coff[994 ] = 64'h000076d0ffffd061;
    assign coff[995 ] = 64'h000076cbffffd056;
    assign coff[996 ] = 64'h000076c7ffffd04a;
    assign coff[997 ] = 64'h000076c2ffffd03e;
    assign coff[998 ] = 64'h000076bdffffd033;
    assign coff[999 ] = 64'h000076b9ffffd027;
    assign coff[1000] = 64'h000076b4ffffd01b;
    assign coff[1001] = 64'h000076afffffd010;
    assign coff[1002] = 64'h000076aaffffd004;
    assign coff[1003] = 64'h000076a6ffffcff8;
    assign coff[1004] = 64'h000076a1ffffcfed;
    assign coff[1005] = 64'h0000769cffffcfe1;
    assign coff[1006] = 64'h00007698ffffcfd6;
    assign coff[1007] = 64'h00007693ffffcfca;
    assign coff[1008] = 64'h0000768effffcfbe;
    assign coff[1009] = 64'h00007689ffffcfb3;
    assign coff[1010] = 64'h00007685ffffcfa7;
    assign coff[1011] = 64'h00007680ffffcf9b;
    assign coff[1012] = 64'h0000767bffffcf90;
    assign coff[1013] = 64'h00007676ffffcf84;
    assign coff[1014] = 64'h00007672ffffcf78;
    assign coff[1015] = 64'h0000766dffffcf6d;
    assign coff[1016] = 64'h00007668ffffcf61;
    assign coff[1017] = 64'h00007663ffffcf56;
    assign coff[1018] = 64'h0000765effffcf4a;
    assign coff[1019] = 64'h0000765affffcf3e;
    assign coff[1020] = 64'h00007655ffffcf33;
    assign coff[1021] = 64'h00007650ffffcf27;
    assign coff[1022] = 64'h0000764bffffcf1b;
    assign coff[1023] = 64'h00007646ffffcf10;
    assign coff[1024] = 64'h00007642ffffcf04;
    assign coff[1025] = 64'h0000763dffffcef9;
    assign coff[1026] = 64'h00007638ffffceed;
    assign coff[1027] = 64'h00007633ffffcee1;
    assign coff[1028] = 64'h0000762effffced6;
    assign coff[1029] = 64'h0000762affffceca;
    assign coff[1030] = 64'h00007625ffffcebf;
    assign coff[1031] = 64'h00007620ffffceb3;
    assign coff[1032] = 64'h0000761bffffcea7;
    assign coff[1033] = 64'h00007616ffffce9c;
    assign coff[1034] = 64'h00007611ffffce90;
    assign coff[1035] = 64'h0000760dffffce85;
    assign coff[1036] = 64'h00007608ffffce79;
    assign coff[1037] = 64'h00007603ffffce6d;
    assign coff[1038] = 64'h000075feffffce62;
    assign coff[1039] = 64'h000075f9ffffce56;
    assign coff[1040] = 64'h000075f4ffffce4b;
    assign coff[1041] = 64'h000075efffffce3f;
    assign coff[1042] = 64'h000075eaffffce34;
    assign coff[1043] = 64'h000075e6ffffce28;
    assign coff[1044] = 64'h000075e1ffffce1c;
    assign coff[1045] = 64'h000075dcffffce11;
    assign coff[1046] = 64'h000075d7ffffce05;
    assign coff[1047] = 64'h000075d2ffffcdfa;
    assign coff[1048] = 64'h000075cdffffcdee;
    assign coff[1049] = 64'h000075c8ffffcde3;
    assign coff[1050] = 64'h000075c3ffffcdd7;
    assign coff[1051] = 64'h000075beffffcdcb;
    assign coff[1052] = 64'h000075b9ffffcdc0;
    assign coff[1053] = 64'h000075b4ffffcdb4;
    assign coff[1054] = 64'h000075afffffcda9;
    assign coff[1055] = 64'h000075aaffffcd9d;
    assign coff[1056] = 64'h000075a6ffffcd92;
    assign coff[1057] = 64'h000075a1ffffcd86;
    assign coff[1058] = 64'h0000759cffffcd7b;
    assign coff[1059] = 64'h00007597ffffcd6f;
    assign coff[1060] = 64'h00007592ffffcd63;
    assign coff[1061] = 64'h0000758dffffcd58;
    assign coff[1062] = 64'h00007588ffffcd4c;
    assign coff[1063] = 64'h00007583ffffcd41;
    assign coff[1064] = 64'h0000757effffcd35;
    assign coff[1065] = 64'h00007579ffffcd2a;
    assign coff[1066] = 64'h00007574ffffcd1e;
    assign coff[1067] = 64'h0000756fffffcd13;
    assign coff[1068] = 64'h0000756affffcd07;
    assign coff[1069] = 64'h00007565ffffccfc;
    assign coff[1070] = 64'h00007560ffffccf0;
    assign coff[1071] = 64'h0000755bffffcce5;
    assign coff[1072] = 64'h00007556ffffccd9;
    assign coff[1073] = 64'h00007551ffffccce;
    assign coff[1074] = 64'h0000754cffffccc2;
    assign coff[1075] = 64'h00007547ffffccb7;
    assign coff[1076] = 64'h00007542ffffccab;
    assign coff[1077] = 64'h0000753dffffcca0;
    assign coff[1078] = 64'h00007538ffffcc94;
    assign coff[1079] = 64'h00007532ffffcc89;
    assign coff[1080] = 64'h0000752dffffcc7d;
    assign coff[1081] = 64'h00007528ffffcc72;
    assign coff[1082] = 64'h00007523ffffcc66;
    assign coff[1083] = 64'h0000751effffcc5b;
    assign coff[1084] = 64'h00007519ffffcc4f;
    assign coff[1085] = 64'h00007514ffffcc44;
    assign coff[1086] = 64'h0000750fffffcc38;
    assign coff[1087] = 64'h0000750affffcc2d;
    assign coff[1088] = 64'h00007505ffffcc21;
    assign coff[1089] = 64'h00007500ffffcc16;
    assign coff[1090] = 64'h000074fbffffcc0a;
    assign coff[1091] = 64'h000074f6ffffcbff;
    assign coff[1092] = 64'h000074f0ffffcbf3;
    assign coff[1093] = 64'h000074ebffffcbe8;
    assign coff[1094] = 64'h000074e6ffffcbdc;
    assign coff[1095] = 64'h000074e1ffffcbd1;
    assign coff[1096] = 64'h000074dcffffcbc5;
    assign coff[1097] = 64'h000074d7ffffcbba;
    assign coff[1098] = 64'h000074d2ffffcbae;
    assign coff[1099] = 64'h000074cdffffcba3;
    assign coff[1100] = 64'h000074c7ffffcb97;
    assign coff[1101] = 64'h000074c2ffffcb8c;
    assign coff[1102] = 64'h000074bdffffcb80;
    assign coff[1103] = 64'h000074b8ffffcb75;
    assign coff[1104] = 64'h000074b3ffffcb69;
    assign coff[1105] = 64'h000074aeffffcb5e;
    assign coff[1106] = 64'h000074a8ffffcb53;
    assign coff[1107] = 64'h000074a3ffffcb47;
    assign coff[1108] = 64'h0000749effffcb3c;
    assign coff[1109] = 64'h00007499ffffcb30;
    assign coff[1110] = 64'h00007494ffffcb25;
    assign coff[1111] = 64'h0000748fffffcb19;
    assign coff[1112] = 64'h00007489ffffcb0e;
    assign coff[1113] = 64'h00007484ffffcb02;
    assign coff[1114] = 64'h0000747fffffcaf7;
    assign coff[1115] = 64'h0000747affffcaec;
    assign coff[1116] = 64'h00007475ffffcae0;
    assign coff[1117] = 64'h0000746fffffcad5;
    assign coff[1118] = 64'h0000746affffcac9;
    assign coff[1119] = 64'h00007465ffffcabe;
    assign coff[1120] = 64'h00007460ffffcab2;
    assign coff[1121] = 64'h0000745affffcaa7;
    assign coff[1122] = 64'h00007455ffffca9c;
    assign coff[1123] = 64'h00007450ffffca90;
    assign coff[1124] = 64'h0000744bffffca85;
    assign coff[1125] = 64'h00007445ffffca79;
    assign coff[1126] = 64'h00007440ffffca6e;
    assign coff[1127] = 64'h0000743bffffca63;
    assign coff[1128] = 64'h00007436ffffca57;
    assign coff[1129] = 64'h00007430ffffca4c;
    assign coff[1130] = 64'h0000742bffffca40;
    assign coff[1131] = 64'h00007426ffffca35;
    assign coff[1132] = 64'h00007421ffffca29;
    assign coff[1133] = 64'h0000741bffffca1e;
    assign coff[1134] = 64'h00007416ffffca13;
    assign coff[1135] = 64'h00007411ffffca07;
    assign coff[1136] = 64'h0000740bffffc9fc;
    assign coff[1137] = 64'h00007406ffffc9f1;
    assign coff[1138] = 64'h00007401ffffc9e5;
    assign coff[1139] = 64'h000073fbffffc9da;
    assign coff[1140] = 64'h000073f6ffffc9ce;
    assign coff[1141] = 64'h000073f1ffffc9c3;
    assign coff[1142] = 64'h000073ebffffc9b8;
    assign coff[1143] = 64'h000073e6ffffc9ac;
    assign coff[1144] = 64'h000073e1ffffc9a1;
    assign coff[1145] = 64'h000073dbffffc995;
    assign coff[1146] = 64'h000073d6ffffc98a;
    assign coff[1147] = 64'h000073d1ffffc97f;
    assign coff[1148] = 64'h000073cbffffc973;
    assign coff[1149] = 64'h000073c6ffffc968;
    assign coff[1150] = 64'h000073c1ffffc95d;
    assign coff[1151] = 64'h000073bbffffc951;
    assign coff[1152] = 64'h000073b6ffffc946;
    assign coff[1153] = 64'h000073b1ffffc93b;
    assign coff[1154] = 64'h000073abffffc92f;
    assign coff[1155] = 64'h000073a6ffffc924;
    assign coff[1156] = 64'h000073a0ffffc918;
    assign coff[1157] = 64'h0000739bffffc90d;
    assign coff[1158] = 64'h00007396ffffc902;
    assign coff[1159] = 64'h00007390ffffc8f6;
    assign coff[1160] = 64'h0000738bffffc8eb;
    assign coff[1161] = 64'h00007385ffffc8e0;
    assign coff[1162] = 64'h00007380ffffc8d4;
    assign coff[1163] = 64'h0000737bffffc8c9;
    assign coff[1164] = 64'h00007375ffffc8be;
    assign coff[1165] = 64'h00007370ffffc8b2;
    assign coff[1166] = 64'h0000736affffc8a7;
    assign coff[1167] = 64'h00007365ffffc89c;
    assign coff[1168] = 64'h0000735fffffc890;
    assign coff[1169] = 64'h0000735affffc885;
    assign coff[1170] = 64'h00007355ffffc87a;
    assign coff[1171] = 64'h0000734fffffc86e;
    assign coff[1172] = 64'h0000734affffc863;
    assign coff[1173] = 64'h00007344ffffc858;
    assign coff[1174] = 64'h0000733fffffc84c;
    assign coff[1175] = 64'h00007339ffffc841;
    assign coff[1176] = 64'h00007334ffffc836;
    assign coff[1177] = 64'h0000732effffc82b;
    assign coff[1178] = 64'h00007329ffffc81f;
    assign coff[1179] = 64'h00007323ffffc814;
    assign coff[1180] = 64'h0000731effffc809;
    assign coff[1181] = 64'h00007318ffffc7fd;
    assign coff[1182] = 64'h00007313ffffc7f2;
    assign coff[1183] = 64'h0000730dffffc7e7;
    assign coff[1184] = 64'h00007308ffffc7db;
    assign coff[1185] = 64'h00007302ffffc7d0;
    assign coff[1186] = 64'h000072fdffffc7c5;
    assign coff[1187] = 64'h000072f7ffffc7ba;
    assign coff[1188] = 64'h000072f2ffffc7ae;
    assign coff[1189] = 64'h000072ecffffc7a3;
    assign coff[1190] = 64'h000072e7ffffc798;
    assign coff[1191] = 64'h000072e1ffffc78c;
    assign coff[1192] = 64'h000072dcffffc781;
    assign coff[1193] = 64'h000072d6ffffc776;
    assign coff[1194] = 64'h000072d0ffffc76b;
    assign coff[1195] = 64'h000072cbffffc75f;
    assign coff[1196] = 64'h000072c5ffffc754;
    assign coff[1197] = 64'h000072c0ffffc749;
    assign coff[1198] = 64'h000072baffffc73e;
    assign coff[1199] = 64'h000072b5ffffc732;
    assign coff[1200] = 64'h000072afffffc727;
    assign coff[1201] = 64'h000072a9ffffc71c;
    assign coff[1202] = 64'h000072a4ffffc710;
    assign coff[1203] = 64'h0000729effffc705;
    assign coff[1204] = 64'h00007299ffffc6fa;
    assign coff[1205] = 64'h00007293ffffc6ef;
    assign coff[1206] = 64'h0000728dffffc6e3;
    assign coff[1207] = 64'h00007288ffffc6d8;
    assign coff[1208] = 64'h00007282ffffc6cd;
    assign coff[1209] = 64'h0000727dffffc6c2;
    assign coff[1210] = 64'h00007277ffffc6b7;
    assign coff[1211] = 64'h00007271ffffc6ab;
    assign coff[1212] = 64'h0000726cffffc6a0;
    assign coff[1213] = 64'h00007266ffffc695;
    assign coff[1214] = 64'h00007260ffffc68a;
    assign coff[1215] = 64'h0000725bffffc67e;
    assign coff[1216] = 64'h00007255ffffc673;
    assign coff[1217] = 64'h00007250ffffc668;
    assign coff[1218] = 64'h0000724affffc65d;
    assign coff[1219] = 64'h00007244ffffc651;
    assign coff[1220] = 64'h0000723fffffc646;
    assign coff[1221] = 64'h00007239ffffc63b;
    assign coff[1222] = 64'h00007233ffffc630;
    assign coff[1223] = 64'h0000722effffc625;
    assign coff[1224] = 64'h00007228ffffc619;
    assign coff[1225] = 64'h00007222ffffc60e;
    assign coff[1226] = 64'h0000721cffffc603;
    assign coff[1227] = 64'h00007217ffffc5f8;
    assign coff[1228] = 64'h00007211ffffc5ed;
    assign coff[1229] = 64'h0000720bffffc5e1;
    assign coff[1230] = 64'h00007206ffffc5d6;
    assign coff[1231] = 64'h00007200ffffc5cb;
    assign coff[1232] = 64'h000071faffffc5c0;
    assign coff[1233] = 64'h000071f5ffffc5b5;
    assign coff[1234] = 64'h000071efffffc5a9;
    assign coff[1235] = 64'h000071e9ffffc59e;
    assign coff[1236] = 64'h000071e3ffffc593;
    assign coff[1237] = 64'h000071deffffc588;
    assign coff[1238] = 64'h000071d8ffffc57d;
    assign coff[1239] = 64'h000071d2ffffc572;
    assign coff[1240] = 64'h000071ccffffc566;
    assign coff[1241] = 64'h000071c7ffffc55b;
    assign coff[1242] = 64'h000071c1ffffc550;
    assign coff[1243] = 64'h000071bbffffc545;
    assign coff[1244] = 64'h000071b5ffffc53a;
    assign coff[1245] = 64'h000071b0ffffc52f;
    assign coff[1246] = 64'h000071aaffffc523;
    assign coff[1247] = 64'h000071a4ffffc518;
    assign coff[1248] = 64'h0000719effffc50d;
    assign coff[1249] = 64'h00007198ffffc502;
    assign coff[1250] = 64'h00007193ffffc4f7;
    assign coff[1251] = 64'h0000718dffffc4ec;
    assign coff[1252] = 64'h00007187ffffc4e0;
    assign coff[1253] = 64'h00007181ffffc4d5;
    assign coff[1254] = 64'h0000717bffffc4ca;
    assign coff[1255] = 64'h00007176ffffc4bf;
    assign coff[1256] = 64'h00007170ffffc4b4;
    assign coff[1257] = 64'h0000716affffc4a9;
    assign coff[1258] = 64'h00007164ffffc49e;
    assign coff[1259] = 64'h0000715effffc493;
    assign coff[1260] = 64'h00007158ffffc487;
    assign coff[1261] = 64'h00007153ffffc47c;
    assign coff[1262] = 64'h0000714dffffc471;
    assign coff[1263] = 64'h00007147ffffc466;
    assign coff[1264] = 64'h00007141ffffc45b;
    assign coff[1265] = 64'h0000713bffffc450;
    assign coff[1266] = 64'h00007135ffffc445;
    assign coff[1267] = 64'h0000712fffffc43a;
    assign coff[1268] = 64'h0000712affffc42e;
    assign coff[1269] = 64'h00007124ffffc423;
    assign coff[1270] = 64'h0000711effffc418;
    assign coff[1271] = 64'h00007118ffffc40d;
    assign coff[1272] = 64'h00007112ffffc402;
    assign coff[1273] = 64'h0000710cffffc3f7;
    assign coff[1274] = 64'h00007106ffffc3ec;
    assign coff[1275] = 64'h00007100ffffc3e1;
    assign coff[1276] = 64'h000070faffffc3d6;
    assign coff[1277] = 64'h000070f5ffffc3cb;
    assign coff[1278] = 64'h000070efffffc3bf;
    assign coff[1279] = 64'h000070e9ffffc3b4;
    assign coff[1280] = 64'h000070e3ffffc3a9;
    assign coff[1281] = 64'h000070ddffffc39e;
    assign coff[1282] = 64'h000070d7ffffc393;
    assign coff[1283] = 64'h000070d1ffffc388;
    assign coff[1284] = 64'h000070cbffffc37d;
    assign coff[1285] = 64'h000070c5ffffc372;
    assign coff[1286] = 64'h000070bfffffc367;
    assign coff[1287] = 64'h000070b9ffffc35c;
    assign coff[1288] = 64'h000070b3ffffc351;
    assign coff[1289] = 64'h000070adffffc346;
    assign coff[1290] = 64'h000070a7ffffc33b;
    assign coff[1291] = 64'h000070a1ffffc330;
    assign coff[1292] = 64'h0000709bffffc324;
    assign coff[1293] = 64'h00007095ffffc319;
    assign coff[1294] = 64'h0000708fffffc30e;
    assign coff[1295] = 64'h00007089ffffc303;
    assign coff[1296] = 64'h00007083ffffc2f8;
    assign coff[1297] = 64'h0000707dffffc2ed;
    assign coff[1298] = 64'h00007077ffffc2e2;
    assign coff[1299] = 64'h00007071ffffc2d7;
    assign coff[1300] = 64'h0000706bffffc2cc;
    assign coff[1301] = 64'h00007065ffffc2c1;
    assign coff[1302] = 64'h0000705fffffc2b6;
    assign coff[1303] = 64'h00007059ffffc2ab;
    assign coff[1304] = 64'h00007053ffffc2a0;
    assign coff[1305] = 64'h0000704dffffc295;
    assign coff[1306] = 64'h00007047ffffc28a;
    assign coff[1307] = 64'h00007041ffffc27f;
    assign coff[1308] = 64'h0000703bffffc274;
    assign coff[1309] = 64'h00007035ffffc269;
    assign coff[1310] = 64'h0000702fffffc25e;
    assign coff[1311] = 64'h00007029ffffc253;
    assign coff[1312] = 64'h00007023ffffc248;
    assign coff[1313] = 64'h0000701dffffc23d;
    assign coff[1314] = 64'h00007017ffffc232;
    assign coff[1315] = 64'h00007011ffffc227;
    assign coff[1316] = 64'h0000700bffffc21c;
    assign coff[1317] = 64'h00007005ffffc211;
    assign coff[1318] = 64'h00006fffffffc206;
    assign coff[1319] = 64'h00006ff9ffffc1fb;
    assign coff[1320] = 64'h00006ff2ffffc1f0;
    assign coff[1321] = 64'h00006fecffffc1e5;
    assign coff[1322] = 64'h00006fe6ffffc1da;
    assign coff[1323] = 64'h00006fe0ffffc1cf;
    assign coff[1324] = 64'h00006fdaffffc1c4;
    assign coff[1325] = 64'h00006fd4ffffc1b9;
    assign coff[1326] = 64'h00006fceffffc1ae;
    assign coff[1327] = 64'h00006fc8ffffc1a3;
    assign coff[1328] = 64'h00006fc2ffffc198;
    assign coff[1329] = 64'h00006fbbffffc18d;
    assign coff[1330] = 64'h00006fb5ffffc182;
    assign coff[1331] = 64'h00006fafffffc177;
    assign coff[1332] = 64'h00006fa9ffffc16c;
    assign coff[1333] = 64'h00006fa3ffffc161;
    assign coff[1334] = 64'h00006f9dffffc156;
    assign coff[1335] = 64'h00006f97ffffc14b;
    assign coff[1336] = 64'h00006f90ffffc140;
    assign coff[1337] = 64'h00006f8affffc135;
    assign coff[1338] = 64'h00006f84ffffc12a;
    assign coff[1339] = 64'h00006f7effffc11f;
    assign coff[1340] = 64'h00006f78ffffc114;
    assign coff[1341] = 64'h00006f72ffffc10a;
    assign coff[1342] = 64'h00006f6bffffc0ff;
    assign coff[1343] = 64'h00006f65ffffc0f4;
    assign coff[1344] = 64'h00006f5fffffc0e9;
    assign coff[1345] = 64'h00006f59ffffc0de;
    assign coff[1346] = 64'h00006f53ffffc0d3;
    assign coff[1347] = 64'h00006f4cffffc0c8;
    assign coff[1348] = 64'h00006f46ffffc0bd;
    assign coff[1349] = 64'h00006f40ffffc0b2;
    assign coff[1350] = 64'h00006f3affffc0a7;
    assign coff[1351] = 64'h00006f34ffffc09c;
    assign coff[1352] = 64'h00006f2dffffc091;
    assign coff[1353] = 64'h00006f27ffffc086;
    assign coff[1354] = 64'h00006f21ffffc07b;
    assign coff[1355] = 64'h00006f1bffffc071;
    assign coff[1356] = 64'h00006f14ffffc066;
    assign coff[1357] = 64'h00006f0effffc05b;
    assign coff[1358] = 64'h00006f08ffffc050;
    assign coff[1359] = 64'h00006f02ffffc045;
    assign coff[1360] = 64'h00006efbffffc03a;
    assign coff[1361] = 64'h00006ef5ffffc02f;
    assign coff[1362] = 64'h00006eefffffc024;
    assign coff[1363] = 64'h00006ee9ffffc019;
    assign coff[1364] = 64'h00006ee2ffffc00f;
    assign coff[1365] = 64'h00006edcffffc004;
    assign coff[1366] = 64'h00006ed6ffffbff9;
    assign coff[1367] = 64'h00006ecfffffbfee;
    assign coff[1368] = 64'h00006ec9ffffbfe3;
    assign coff[1369] = 64'h00006ec3ffffbfd8;
    assign coff[1370] = 64'h00006ebdffffbfcd;
    assign coff[1371] = 64'h00006eb6ffffbfc2;
    assign coff[1372] = 64'h00006eb0ffffbfb8;
    assign coff[1373] = 64'h00006eaaffffbfad;
    assign coff[1374] = 64'h00006ea3ffffbfa2;
    assign coff[1375] = 64'h00006e9dffffbf97;
    assign coff[1376] = 64'h00006e97ffffbf8c;
    assign coff[1377] = 64'h00006e90ffffbf81;
    assign coff[1378] = 64'h00006e8affffbf76;
    assign coff[1379] = 64'h00006e84ffffbf6b;
    assign coff[1380] = 64'h00006e7dffffbf61;
    assign coff[1381] = 64'h00006e77ffffbf56;
    assign coff[1382] = 64'h00006e71ffffbf4b;
    assign coff[1383] = 64'h00006e6affffbf40;
    assign coff[1384] = 64'h00006e64ffffbf35;
    assign coff[1385] = 64'h00006e5effffbf2a;
    assign coff[1386] = 64'h00006e57ffffbf20;
    assign coff[1387] = 64'h00006e51ffffbf15;
    assign coff[1388] = 64'h00006e4affffbf0a;
    assign coff[1389] = 64'h00006e44ffffbeff;
    assign coff[1390] = 64'h00006e3effffbef4;
    assign coff[1391] = 64'h00006e37ffffbee9;
    assign coff[1392] = 64'h00006e31ffffbedf;
    assign coff[1393] = 64'h00006e2affffbed4;
    assign coff[1394] = 64'h00006e24ffffbec9;
    assign coff[1395] = 64'h00006e1effffbebe;
    assign coff[1396] = 64'h00006e17ffffbeb3;
    assign coff[1397] = 64'h00006e11ffffbea9;
    assign coff[1398] = 64'h00006e0affffbe9e;
    assign coff[1399] = 64'h00006e04ffffbe93;
    assign coff[1400] = 64'h00006dfeffffbe88;
    assign coff[1401] = 64'h00006df7ffffbe7d;
    assign coff[1402] = 64'h00006df1ffffbe73;
    assign coff[1403] = 64'h00006deaffffbe68;
    assign coff[1404] = 64'h00006de4ffffbe5d;
    assign coff[1405] = 64'h00006dddffffbe52;
    assign coff[1406] = 64'h00006dd7ffffbe47;
    assign coff[1407] = 64'h00006dd1ffffbe3d;
    assign coff[1408] = 64'h00006dcaffffbe32;
    assign coff[1409] = 64'h00006dc4ffffbe27;
    assign coff[1410] = 64'h00006dbdffffbe1c;
    assign coff[1411] = 64'h00006db7ffffbe12;
    assign coff[1412] = 64'h00006db0ffffbe07;
    assign coff[1413] = 64'h00006daaffffbdfc;
    assign coff[1414] = 64'h00006da3ffffbdf1;
    assign coff[1415] = 64'h00006d9dffffbde6;
    assign coff[1416] = 64'h00006d96ffffbddc;
    assign coff[1417] = 64'h00006d90ffffbdd1;
    assign coff[1418] = 64'h00006d89ffffbdc6;
    assign coff[1419] = 64'h00006d83ffffbdbb;
    assign coff[1420] = 64'h00006d7cffffbdb1;
    assign coff[1421] = 64'h00006d76ffffbda6;
    assign coff[1422] = 64'h00006d6fffffbd9b;
    assign coff[1423] = 64'h00006d69ffffbd90;
    assign coff[1424] = 64'h00006d62ffffbd86;
    assign coff[1425] = 64'h00006d5cffffbd7b;
    assign coff[1426] = 64'h00006d55ffffbd70;
    assign coff[1427] = 64'h00006d4fffffbd66;
    assign coff[1428] = 64'h00006d48ffffbd5b;
    assign coff[1429] = 64'h00006d41ffffbd50;
    assign coff[1430] = 64'h00006d3bffffbd45;
    assign coff[1431] = 64'h00006d34ffffbd3b;
    assign coff[1432] = 64'h00006d2effffbd30;
    assign coff[1433] = 64'h00006d27ffffbd25;
    assign coff[1434] = 64'h00006d21ffffbd1a;
    assign coff[1435] = 64'h00006d1affffbd10;
    assign coff[1436] = 64'h00006d14ffffbd05;
    assign coff[1437] = 64'h00006d0dffffbcfa;
    assign coff[1438] = 64'h00006d06ffffbcf0;
    assign coff[1439] = 64'h00006d00ffffbce5;
    assign coff[1440] = 64'h00006cf9ffffbcda;
    assign coff[1441] = 64'h00006cf3ffffbcd0;
    assign coff[1442] = 64'h00006cecffffbcc5;
    assign coff[1443] = 64'h00006ce5ffffbcba;
    assign coff[1444] = 64'h00006cdfffffbcaf;
    assign coff[1445] = 64'h00006cd8ffffbca5;
    assign coff[1446] = 64'h00006cd2ffffbc9a;
    assign coff[1447] = 64'h00006ccbffffbc8f;
    assign coff[1448] = 64'h00006cc4ffffbc85;
    assign coff[1449] = 64'h00006cbeffffbc7a;
    assign coff[1450] = 64'h00006cb7ffffbc6f;
    assign coff[1451] = 64'h00006cb0ffffbc65;
    assign coff[1452] = 64'h00006caaffffbc5a;
    assign coff[1453] = 64'h00006ca3ffffbc4f;
    assign coff[1454] = 64'h00006c9dffffbc45;
    assign coff[1455] = 64'h00006c96ffffbc3a;
    assign coff[1456] = 64'h00006c8fffffbc2f;
    assign coff[1457] = 64'h00006c89ffffbc25;
    assign coff[1458] = 64'h00006c82ffffbc1a;
    assign coff[1459] = 64'h00006c7bffffbc0f;
    assign coff[1460] = 64'h00006c75ffffbc05;
    assign coff[1461] = 64'h00006c6effffbbfa;
    assign coff[1462] = 64'h00006c67ffffbbef;
    assign coff[1463] = 64'h00006c61ffffbbe5;
    assign coff[1464] = 64'h00006c5affffbbda;
    assign coff[1465] = 64'h00006c53ffffbbd0;
    assign coff[1466] = 64'h00006c4cffffbbc5;
    assign coff[1467] = 64'h00006c46ffffbbba;
    assign coff[1468] = 64'h00006c3fffffbbb0;
    assign coff[1469] = 64'h00006c38ffffbba5;
    assign coff[1470] = 64'h00006c32ffffbb9a;
    assign coff[1471] = 64'h00006c2bffffbb90;
    assign coff[1472] = 64'h00006c24ffffbb85;
    assign coff[1473] = 64'h00006c1dffffbb7b;
    assign coff[1474] = 64'h00006c17ffffbb70;
    assign coff[1475] = 64'h00006c10ffffbb65;
    assign coff[1476] = 64'h00006c09ffffbb5b;
    assign coff[1477] = 64'h00006c02ffffbb50;
    assign coff[1478] = 64'h00006bfcffffbb46;
    assign coff[1479] = 64'h00006bf5ffffbb3b;
    assign coff[1480] = 64'h00006beeffffbb30;
    assign coff[1481] = 64'h00006be7ffffbb26;
    assign coff[1482] = 64'h00006be1ffffbb1b;
    assign coff[1483] = 64'h00006bdaffffbb11;
    assign coff[1484] = 64'h00006bd3ffffbb06;
    assign coff[1485] = 64'h00006bccffffbafb;
    assign coff[1486] = 64'h00006bc6ffffbaf1;
    assign coff[1487] = 64'h00006bbfffffbae6;
    assign coff[1488] = 64'h00006bb8ffffbadc;
    assign coff[1489] = 64'h00006bb1ffffbad1;
    assign coff[1490] = 64'h00006baaffffbac7;
    assign coff[1491] = 64'h00006ba4ffffbabc;
    assign coff[1492] = 64'h00006b9dffffbab1;
    assign coff[1493] = 64'h00006b96ffffbaa7;
    assign coff[1494] = 64'h00006b8fffffba9c;
    assign coff[1495] = 64'h00006b88ffffba92;
    assign coff[1496] = 64'h00006b82ffffba87;
    assign coff[1497] = 64'h00006b7bffffba7d;
    assign coff[1498] = 64'h00006b74ffffba72;
    assign coff[1499] = 64'h00006b6dffffba67;
    assign coff[1500] = 64'h00006b66ffffba5d;
    assign coff[1501] = 64'h00006b5fffffba52;
    assign coff[1502] = 64'h00006b59ffffba48;
    assign coff[1503] = 64'h00006b52ffffba3d;
    assign coff[1504] = 64'h00006b4bffffba33;
    assign coff[1505] = 64'h00006b44ffffba28;
    assign coff[1506] = 64'h00006b3dffffba1e;
    assign coff[1507] = 64'h00006b36ffffba13;
    assign coff[1508] = 64'h00006b30ffffba09;
    assign coff[1509] = 64'h00006b29ffffb9fe;
    assign coff[1510] = 64'h00006b22ffffb9f4;
    assign coff[1511] = 64'h00006b1bffffb9e9;
    assign coff[1512] = 64'h00006b14ffffb9df;
    assign coff[1513] = 64'h00006b0dffffb9d4;
    assign coff[1514] = 64'h00006b06ffffb9ca;
    assign coff[1515] = 64'h00006affffffb9bf;
    assign coff[1516] = 64'h00006af8ffffb9b5;
    assign coff[1517] = 64'h00006af2ffffb9aa;
    assign coff[1518] = 64'h00006aebffffb9a0;
    assign coff[1519] = 64'h00006ae4ffffb995;
    assign coff[1520] = 64'h00006addffffb98b;
    assign coff[1521] = 64'h00006ad6ffffb980;
    assign coff[1522] = 64'h00006acfffffb976;
    assign coff[1523] = 64'h00006ac8ffffb96b;
    assign coff[1524] = 64'h00006ac1ffffb961;
    assign coff[1525] = 64'h00006abaffffb956;
    assign coff[1526] = 64'h00006ab3ffffb94c;
    assign coff[1527] = 64'h00006aacffffb941;
    assign coff[1528] = 64'h00006aa5ffffb937;
    assign coff[1529] = 64'h00006a9effffb92c;
    assign coff[1530] = 64'h00006a97ffffb922;
    assign coff[1531] = 64'h00006a90ffffb917;
    assign coff[1532] = 64'h00006a89ffffb90d;
    assign coff[1533] = 64'h00006a83ffffb902;
    assign coff[1534] = 64'h00006a7cffffb8f8;
    assign coff[1535] = 64'h00006a75ffffb8ee;
    assign coff[1536] = 64'h00006a6effffb8e3;
    assign coff[1537] = 64'h00006a67ffffb8d9;
    assign coff[1538] = 64'h00006a60ffffb8ce;
    assign coff[1539] = 64'h00006a59ffffb8c4;
    assign coff[1540] = 64'h00006a52ffffb8b9;
    assign coff[1541] = 64'h00006a4bffffb8af;
    assign coff[1542] = 64'h00006a44ffffb8a4;
    assign coff[1543] = 64'h00006a3dffffb89a;
    assign coff[1544] = 64'h00006a36ffffb890;
    assign coff[1545] = 64'h00006a2fffffb885;
    assign coff[1546] = 64'h00006a28ffffb87b;
    assign coff[1547] = 64'h00006a21ffffb870;
    assign coff[1548] = 64'h00006a1affffb866;
    assign coff[1549] = 64'h00006a12ffffb85b;
    assign coff[1550] = 64'h00006a0bffffb851;
    assign coff[1551] = 64'h00006a04ffffb847;
    assign coff[1552] = 64'h000069fdffffb83c;
    assign coff[1553] = 64'h000069f6ffffb832;
    assign coff[1554] = 64'h000069efffffb827;
    assign coff[1555] = 64'h000069e8ffffb81d;
    assign coff[1556] = 64'h000069e1ffffb813;
    assign coff[1557] = 64'h000069daffffb808;
    assign coff[1558] = 64'h000069d3ffffb7fe;
    assign coff[1559] = 64'h000069ccffffb7f3;
    assign coff[1560] = 64'h000069c5ffffb7e9;
    assign coff[1561] = 64'h000069beffffb7df;
    assign coff[1562] = 64'h000069b7ffffb7d4;
    assign coff[1563] = 64'h000069b0ffffb7ca;
    assign coff[1564] = 64'h000069a9ffffb7c0;
    assign coff[1565] = 64'h000069a1ffffb7b5;
    assign coff[1566] = 64'h0000699affffb7ab;
    assign coff[1567] = 64'h00006993ffffb7a0;
    assign coff[1568] = 64'h0000698cffffb796;
    assign coff[1569] = 64'h00006985ffffb78c;
    assign coff[1570] = 64'h0000697effffb781;
    assign coff[1571] = 64'h00006977ffffb777;
    assign coff[1572] = 64'h00006970ffffb76d;
    assign coff[1573] = 64'h00006969ffffb762;
    assign coff[1574] = 64'h00006961ffffb758;
    assign coff[1575] = 64'h0000695affffb74e;
    assign coff[1576] = 64'h00006953ffffb743;
    assign coff[1577] = 64'h0000694cffffb739;
    assign coff[1578] = 64'h00006945ffffb72f;
    assign coff[1579] = 64'h0000693effffb724;
    assign coff[1580] = 64'h00006937ffffb71a;
    assign coff[1581] = 64'h0000692fffffb710;
    assign coff[1582] = 64'h00006928ffffb705;
    assign coff[1583] = 64'h00006921ffffb6fb;
    assign coff[1584] = 64'h0000691affffb6f1;
    assign coff[1585] = 64'h00006913ffffb6e6;
    assign coff[1586] = 64'h0000690cffffb6dc;
    assign coff[1587] = 64'h00006904ffffb6d2;
    assign coff[1588] = 64'h000068fdffffb6c7;
    assign coff[1589] = 64'h000068f6ffffb6bd;
    assign coff[1590] = 64'h000068efffffb6b3;
    assign coff[1591] = 64'h000068e8ffffb6a8;
    assign coff[1592] = 64'h000068e0ffffb69e;
    assign coff[1593] = 64'h000068d9ffffb694;
    assign coff[1594] = 64'h000068d2ffffb68a;
    assign coff[1595] = 64'h000068cbffffb67f;
    assign coff[1596] = 64'h000068c4ffffb675;
    assign coff[1597] = 64'h000068bcffffb66b;
    assign coff[1598] = 64'h000068b5ffffb660;
    assign coff[1599] = 64'h000068aeffffb656;
    assign coff[1600] = 64'h000068a7ffffb64c;
    assign coff[1601] = 64'h0000689fffffb642;
    assign coff[1602] = 64'h00006898ffffb637;
    assign coff[1603] = 64'h00006891ffffb62d;
    assign coff[1604] = 64'h0000688affffb623;
    assign coff[1605] = 64'h00006882ffffb619;
    assign coff[1606] = 64'h0000687bffffb60e;
    assign coff[1607] = 64'h00006874ffffb604;
    assign coff[1608] = 64'h0000686dffffb5fa;
    assign coff[1609] = 64'h00006865ffffb5f0;
    assign coff[1610] = 64'h0000685effffb5e5;
    assign coff[1611] = 64'h00006857ffffb5db;
    assign coff[1612] = 64'h00006850ffffb5d1;
    assign coff[1613] = 64'h00006848ffffb5c7;
    assign coff[1614] = 64'h00006841ffffb5bc;
    assign coff[1615] = 64'h0000683affffb5b2;
    assign coff[1616] = 64'h00006832ffffb5a8;
    assign coff[1617] = 64'h0000682bffffb59e;
    assign coff[1618] = 64'h00006824ffffb593;
    assign coff[1619] = 64'h0000681cffffb589;
    assign coff[1620] = 64'h00006815ffffb57f;
    assign coff[1621] = 64'h0000680effffb575;
    assign coff[1622] = 64'h00006806ffffb56b;
    assign coff[1623] = 64'h000067ffffffb560;
    assign coff[1624] = 64'h000067f8ffffb556;
    assign coff[1625] = 64'h000067f0ffffb54c;
    assign coff[1626] = 64'h000067e9ffffb542;
    assign coff[1627] = 64'h000067e2ffffb538;
    assign coff[1628] = 64'h000067daffffb52d;
    assign coff[1629] = 64'h000067d3ffffb523;
    assign coff[1630] = 64'h000067ccffffb519;
    assign coff[1631] = 64'h000067c4ffffb50f;
    assign coff[1632] = 64'h000067bdffffb505;
    assign coff[1633] = 64'h000067b6ffffb4fa;
    assign coff[1634] = 64'h000067aeffffb4f0;
    assign coff[1635] = 64'h000067a7ffffb4e6;
    assign coff[1636] = 64'h000067a0ffffb4dc;
    assign coff[1637] = 64'h00006798ffffb4d2;
    assign coff[1638] = 64'h00006791ffffb4c8;
    assign coff[1639] = 64'h00006789ffffb4bd;
    assign coff[1640] = 64'h00006782ffffb4b3;
    assign coff[1641] = 64'h0000677bffffb4a9;
    assign coff[1642] = 64'h00006773ffffb49f;
    assign coff[1643] = 64'h0000676cffffb495;
    assign coff[1644] = 64'h00006764ffffb48b;
    assign coff[1645] = 64'h0000675dffffb480;
    assign coff[1646] = 64'h00006756ffffb476;
    assign coff[1647] = 64'h0000674effffb46c;
    assign coff[1648] = 64'h00006747ffffb462;
    assign coff[1649] = 64'h0000673fffffb458;
    assign coff[1650] = 64'h00006738ffffb44e;
    assign coff[1651] = 64'h00006730ffffb444;
    assign coff[1652] = 64'h00006729ffffb439;
    assign coff[1653] = 64'h00006722ffffb42f;
    assign coff[1654] = 64'h0000671affffb425;
    assign coff[1655] = 64'h00006713ffffb41b;
    assign coff[1656] = 64'h0000670bffffb411;
    assign coff[1657] = 64'h00006704ffffb407;
    assign coff[1658] = 64'h000066fcffffb3fd;
    assign coff[1659] = 64'h000066f5ffffb3f3;
    assign coff[1660] = 64'h000066edffffb3e9;
    assign coff[1661] = 64'h000066e6ffffb3de;
    assign coff[1662] = 64'h000066deffffb3d4;
    assign coff[1663] = 64'h000066d7ffffb3ca;
    assign coff[1664] = 64'h000066d0ffffb3c0;
    assign coff[1665] = 64'h000066c8ffffb3b6;
    assign coff[1666] = 64'h000066c1ffffb3ac;
    assign coff[1667] = 64'h000066b9ffffb3a2;
    assign coff[1668] = 64'h000066b2ffffb398;
    assign coff[1669] = 64'h000066aaffffb38e;
    assign coff[1670] = 64'h000066a3ffffb384;
    assign coff[1671] = 64'h0000669bffffb37a;
    assign coff[1672] = 64'h00006693ffffb36f;
    assign coff[1673] = 64'h0000668cffffb365;
    assign coff[1674] = 64'h00006684ffffb35b;
    assign coff[1675] = 64'h0000667dffffb351;
    assign coff[1676] = 64'h00006675ffffb347;
    assign coff[1677] = 64'h0000666effffb33d;
    assign coff[1678] = 64'h00006666ffffb333;
    assign coff[1679] = 64'h0000665fffffb329;
    assign coff[1680] = 64'h00006657ffffb31f;
    assign coff[1681] = 64'h00006650ffffb315;
    assign coff[1682] = 64'h00006648ffffb30b;
    assign coff[1683] = 64'h00006641ffffb301;
    assign coff[1684] = 64'h00006639ffffb2f7;
    assign coff[1685] = 64'h00006631ffffb2ed;
    assign coff[1686] = 64'h0000662affffb2e3;
    assign coff[1687] = 64'h00006622ffffb2d9;
    assign coff[1688] = 64'h0000661bffffb2cf;
    assign coff[1689] = 64'h00006613ffffb2c5;
    assign coff[1690] = 64'h0000660cffffb2bb;
    assign coff[1691] = 64'h00006604ffffb2b1;
    assign coff[1692] = 64'h000065fcffffb2a7;
    assign coff[1693] = 64'h000065f5ffffb29d;
    assign coff[1694] = 64'h000065edffffb293;
    assign coff[1695] = 64'h000065e6ffffb289;
    assign coff[1696] = 64'h000065deffffb27f;
    assign coff[1697] = 64'h000065d6ffffb275;
    assign coff[1698] = 64'h000065cfffffb26b;
    assign coff[1699] = 64'h000065c7ffffb261;
    assign coff[1700] = 64'h000065c0ffffb257;
    assign coff[1701] = 64'h000065b8ffffb24d;
    assign coff[1702] = 64'h000065b0ffffb243;
    assign coff[1703] = 64'h000065a9ffffb239;
    assign coff[1704] = 64'h000065a1ffffb22f;
    assign coff[1705] = 64'h00006599ffffb225;
    assign coff[1706] = 64'h00006592ffffb21b;
    assign coff[1707] = 64'h0000658affffb211;
    assign coff[1708] = 64'h00006582ffffb207;
    assign coff[1709] = 64'h0000657bffffb1fd;
    assign coff[1710] = 64'h00006573ffffb1f3;
    assign coff[1711] = 64'h0000656bffffb1e9;
    assign coff[1712] = 64'h00006564ffffb1df;
    assign coff[1713] = 64'h0000655cffffb1d5;
    assign coff[1714] = 64'h00006554ffffb1cb;
    assign coff[1715] = 64'h0000654dffffb1c1;
    assign coff[1716] = 64'h00006545ffffb1b7;
    assign coff[1717] = 64'h0000653dffffb1ad;
    assign coff[1718] = 64'h00006536ffffb1a3;
    assign coff[1719] = 64'h0000652effffb199;
    assign coff[1720] = 64'h00006526ffffb18f;
    assign coff[1721] = 64'h0000651fffffb186;
    assign coff[1722] = 64'h00006517ffffb17c;
    assign coff[1723] = 64'h0000650fffffb172;
    assign coff[1724] = 64'h00006507ffffb168;
    assign coff[1725] = 64'h00006500ffffb15e;
    assign coff[1726] = 64'h000064f8ffffb154;
    assign coff[1727] = 64'h000064f0ffffb14a;
    assign coff[1728] = 64'h000064e9ffffb140;
    assign coff[1729] = 64'h000064e1ffffb136;
    assign coff[1730] = 64'h000064d9ffffb12c;
    assign coff[1731] = 64'h000064d1ffffb122;
    assign coff[1732] = 64'h000064caffffb118;
    assign coff[1733] = 64'h000064c2ffffb10f;
    assign coff[1734] = 64'h000064baffffb105;
    assign coff[1735] = 64'h000064b2ffffb0fb;
    assign coff[1736] = 64'h000064abffffb0f1;
    assign coff[1737] = 64'h000064a3ffffb0e7;
    assign coff[1738] = 64'h0000649bffffb0dd;
    assign coff[1739] = 64'h00006493ffffb0d3;
    assign coff[1740] = 64'h0000648bffffb0c9;
    assign coff[1741] = 64'h00006484ffffb0c0;
    assign coff[1742] = 64'h0000647cffffb0b6;
    assign coff[1743] = 64'h00006474ffffb0ac;
    assign coff[1744] = 64'h0000646cffffb0a2;
    assign coff[1745] = 64'h00006465ffffb098;
    assign coff[1746] = 64'h0000645dffffb08e;
    assign coff[1747] = 64'h00006455ffffb084;
    assign coff[1748] = 64'h0000644dffffb07b;
    assign coff[1749] = 64'h00006445ffffb071;
    assign coff[1750] = 64'h0000643effffb067;
    assign coff[1751] = 64'h00006436ffffb05d;
    assign coff[1752] = 64'h0000642effffb053;
    assign coff[1753] = 64'h00006426ffffb049;
    assign coff[1754] = 64'h0000641effffb040;
    assign coff[1755] = 64'h00006416ffffb036;
    assign coff[1756] = 64'h0000640fffffb02c;
    assign coff[1757] = 64'h00006407ffffb022;
    assign coff[1758] = 64'h000063ffffffb018;
    assign coff[1759] = 64'h000063f7ffffb00e;
    assign coff[1760] = 64'h000063efffffb005;
    assign coff[1761] = 64'h000063e7ffffaffb;
    assign coff[1762] = 64'h000063dfffffaff1;
    assign coff[1763] = 64'h000063d8ffffafe7;
    assign coff[1764] = 64'h000063d0ffffafdd;
    assign coff[1765] = 64'h000063c8ffffafd4;
    assign coff[1766] = 64'h000063c0ffffafca;
    assign coff[1767] = 64'h000063b8ffffafc0;
    assign coff[1768] = 64'h000063b0ffffafb6;
    assign coff[1769] = 64'h000063a8ffffafac;
    assign coff[1770] = 64'h000063a0ffffafa3;
    assign coff[1771] = 64'h00006399ffffaf99;
    assign coff[1772] = 64'h00006391ffffaf8f;
    assign coff[1773] = 64'h00006389ffffaf85;
    assign coff[1774] = 64'h00006381ffffaf7c;
    assign coff[1775] = 64'h00006379ffffaf72;
    assign coff[1776] = 64'h00006371ffffaf68;
    assign coff[1777] = 64'h00006369ffffaf5e;
    assign coff[1778] = 64'h00006361ffffaf54;
    assign coff[1779] = 64'h00006359ffffaf4b;
    assign coff[1780] = 64'h00006351ffffaf41;
    assign coff[1781] = 64'h00006349ffffaf37;
    assign coff[1782] = 64'h00006342ffffaf2d;
    assign coff[1783] = 64'h0000633affffaf24;
    assign coff[1784] = 64'h00006332ffffaf1a;
    assign coff[1785] = 64'h0000632affffaf10;
    assign coff[1786] = 64'h00006322ffffaf07;
    assign coff[1787] = 64'h0000631affffaefd;
    assign coff[1788] = 64'h00006312ffffaef3;
    assign coff[1789] = 64'h0000630affffaee9;
    assign coff[1790] = 64'h00006302ffffaee0;
    assign coff[1791] = 64'h000062faffffaed6;
    assign coff[1792] = 64'h000062f2ffffaecc;
    assign coff[1793] = 64'h000062eaffffaec2;
    assign coff[1794] = 64'h000062e2ffffaeb9;
    assign coff[1795] = 64'h000062daffffaeaf;
    assign coff[1796] = 64'h000062d2ffffaea5;
    assign coff[1797] = 64'h000062caffffae9c;
    assign coff[1798] = 64'h000062c2ffffae92;
    assign coff[1799] = 64'h000062baffffae88;
    assign coff[1800] = 64'h000062b2ffffae7f;
    assign coff[1801] = 64'h000062aaffffae75;
    assign coff[1802] = 64'h000062a2ffffae6b;
    assign coff[1803] = 64'h0000629affffae62;
    assign coff[1804] = 64'h00006292ffffae58;
    assign coff[1805] = 64'h0000628affffae4e;
    assign coff[1806] = 64'h00006282ffffae45;
    assign coff[1807] = 64'h0000627affffae3b;
    assign coff[1808] = 64'h00006272ffffae31;
    assign coff[1809] = 64'h0000626affffae28;
    assign coff[1810] = 64'h00006262ffffae1e;
    assign coff[1811] = 64'h0000625affffae14;
    assign coff[1812] = 64'h00006252ffffae0b;
    assign coff[1813] = 64'h0000624affffae01;
    assign coff[1814] = 64'h00006242ffffadf7;
    assign coff[1815] = 64'h0000623affffadee;
    assign coff[1816] = 64'h00006232ffffade4;
    assign coff[1817] = 64'h0000622affffadda;
    assign coff[1818] = 64'h00006221ffffadd1;
    assign coff[1819] = 64'h00006219ffffadc7;
    assign coff[1820] = 64'h00006211ffffadbd;
    assign coff[1821] = 64'h00006209ffffadb4;
    assign coff[1822] = 64'h00006201ffffadaa;
    assign coff[1823] = 64'h000061f9ffffada1;
    assign coff[1824] = 64'h000061f1ffffad97;
    assign coff[1825] = 64'h000061e9ffffad8d;
    assign coff[1826] = 64'h000061e1ffffad84;
    assign coff[1827] = 64'h000061d9ffffad7a;
    assign coff[1828] = 64'h000061d1ffffad70;
    assign coff[1829] = 64'h000061c9ffffad67;
    assign coff[1830] = 64'h000061c0ffffad5d;
    assign coff[1831] = 64'h000061b8ffffad54;
    assign coff[1832] = 64'h000061b0ffffad4a;
    assign coff[1833] = 64'h000061a8ffffad41;
    assign coff[1834] = 64'h000061a0ffffad37;
    assign coff[1835] = 64'h00006198ffffad2d;
    assign coff[1836] = 64'h00006190ffffad24;
    assign coff[1837] = 64'h00006188ffffad1a;
    assign coff[1838] = 64'h0000617fffffad11;
    assign coff[1839] = 64'h00006177ffffad07;
    assign coff[1840] = 64'h0000616fffffacfd;
    assign coff[1841] = 64'h00006167ffffacf4;
    assign coff[1842] = 64'h0000615fffffacea;
    assign coff[1843] = 64'h00006157fffface1;
    assign coff[1844] = 64'h0000614effffacd7;
    assign coff[1845] = 64'h00006146ffffacce;
    assign coff[1846] = 64'h0000613effffacc4;
    assign coff[1847] = 64'h00006136ffffacbb;
    assign coff[1848] = 64'h0000612effffacb1;
    assign coff[1849] = 64'h00006126ffffaca8;
    assign coff[1850] = 64'h0000611dffffac9e;
    assign coff[1851] = 64'h00006115ffffac94;
    assign coff[1852] = 64'h0000610dffffac8b;
    assign coff[1853] = 64'h00006105ffffac81;
    assign coff[1854] = 64'h000060fdffffac78;
    assign coff[1855] = 64'h000060f4ffffac6e;
    assign coff[1856] = 64'h000060ecffffac65;
    assign coff[1857] = 64'h000060e4ffffac5b;
    assign coff[1858] = 64'h000060dcffffac52;
    assign coff[1859] = 64'h000060d4ffffac48;
    assign coff[1860] = 64'h000060cbffffac3f;
    assign coff[1861] = 64'h000060c3ffffac35;
    assign coff[1862] = 64'h000060bbffffac2c;
    assign coff[1863] = 64'h000060b3ffffac22;
    assign coff[1864] = 64'h000060aaffffac19;
    assign coff[1865] = 64'h000060a2ffffac0f;
    assign coff[1866] = 64'h0000609affffac06;
    assign coff[1867] = 64'h00006092ffffabfc;
    assign coff[1868] = 64'h00006089ffffabf3;
    assign coff[1869] = 64'h00006081ffffabe9;
    assign coff[1870] = 64'h00006079ffffabe0;
    assign coff[1871] = 64'h00006071ffffabd6;
    assign coff[1872] = 64'h00006068ffffabcd;
    assign coff[1873] = 64'h00006060ffffabc4;
    assign coff[1874] = 64'h00006058ffffabba;
    assign coff[1875] = 64'h00006050ffffabb1;
    assign coff[1876] = 64'h00006047ffffaba7;
    assign coff[1877] = 64'h0000603fffffab9e;
    assign coff[1878] = 64'h00006037ffffab94;
    assign coff[1879] = 64'h0000602effffab8b;
    assign coff[1880] = 64'h00006026ffffab81;
    assign coff[1881] = 64'h0000601effffab78;
    assign coff[1882] = 64'h00006016ffffab6f;
    assign coff[1883] = 64'h0000600dffffab65;
    assign coff[1884] = 64'h00006005ffffab5c;
    assign coff[1885] = 64'h00005ffdffffab52;
    assign coff[1886] = 64'h00005ff4ffffab49;
    assign coff[1887] = 64'h00005fecffffab3f;
    assign coff[1888] = 64'h00005fe4ffffab36;
    assign coff[1889] = 64'h00005fdbffffab2d;
    assign coff[1890] = 64'h00005fd3ffffab23;
    assign coff[1891] = 64'h00005fcbffffab1a;
    assign coff[1892] = 64'h00005fc2ffffab10;
    assign coff[1893] = 64'h00005fbaffffab07;
    assign coff[1894] = 64'h00005fb2ffffaafe;
    assign coff[1895] = 64'h00005fa9ffffaaf4;
    assign coff[1896] = 64'h00005fa1ffffaaeb;
    assign coff[1897] = 64'h00005f99ffffaae1;
    assign coff[1898] = 64'h00005f90ffffaad8;
    assign coff[1899] = 64'h00005f88ffffaacf;
    assign coff[1900] = 64'h00005f80ffffaac5;
    assign coff[1901] = 64'h00005f77ffffaabc;
    assign coff[1902] = 64'h00005f6fffffaab2;
    assign coff[1903] = 64'h00005f66ffffaaa9;
    assign coff[1904] = 64'h00005f5effffaaa0;
    assign coff[1905] = 64'h00005f56ffffaa96;
    assign coff[1906] = 64'h00005f4dffffaa8d;
    assign coff[1907] = 64'h00005f45ffffaa84;
    assign coff[1908] = 64'h00005f3cffffaa7a;
    assign coff[1909] = 64'h00005f34ffffaa71;
    assign coff[1910] = 64'h00005f2cffffaa68;
    assign coff[1911] = 64'h00005f23ffffaa5e;
    assign coff[1912] = 64'h00005f1bffffaa55;
    assign coff[1913] = 64'h00005f12ffffaa4c;
    assign coff[1914] = 64'h00005f0affffaa42;
    assign coff[1915] = 64'h00005f02ffffaa39;
    assign coff[1916] = 64'h00005ef9ffffaa30;
    assign coff[1917] = 64'h00005ef1ffffaa26;
    assign coff[1918] = 64'h00005ee8ffffaa1d;
    assign coff[1919] = 64'h00005ee0ffffaa14;
    assign coff[1920] = 64'h00005ed7ffffaa0a;
    assign coff[1921] = 64'h00005ecfffffaa01;
    assign coff[1922] = 64'h00005ec7ffffa9f8;
    assign coff[1923] = 64'h00005ebeffffa9ee;
    assign coff[1924] = 64'h00005eb6ffffa9e5;
    assign coff[1925] = 64'h00005eadffffa9dc;
    assign coff[1926] = 64'h00005ea5ffffa9d3;
    assign coff[1927] = 64'h00005e9cffffa9c9;
    assign coff[1928] = 64'h00005e94ffffa9c0;
    assign coff[1929] = 64'h00005e8bffffa9b7;
    assign coff[1930] = 64'h00005e83ffffa9ad;
    assign coff[1931] = 64'h00005e7affffa9a4;
    assign coff[1932] = 64'h00005e72ffffa99b;
    assign coff[1933] = 64'h00005e69ffffa992;
    assign coff[1934] = 64'h00005e61ffffa988;
    assign coff[1935] = 64'h00005e58ffffa97f;
    assign coff[1936] = 64'h00005e50ffffa976;
    assign coff[1937] = 64'h00005e48ffffa96d;
    assign coff[1938] = 64'h00005e3fffffa963;
    assign coff[1939] = 64'h00005e37ffffa95a;
    assign coff[1940] = 64'h00005e2effffa951;
    assign coff[1941] = 64'h00005e25ffffa948;
    assign coff[1942] = 64'h00005e1dffffa93e;
    assign coff[1943] = 64'h00005e14ffffa935;
    assign coff[1944] = 64'h00005e0cffffa92c;
    assign coff[1945] = 64'h00005e03ffffa923;
    assign coff[1946] = 64'h00005dfbffffa919;
    assign coff[1947] = 64'h00005df2ffffa910;
    assign coff[1948] = 64'h00005deaffffa907;
    assign coff[1949] = 64'h00005de1ffffa8fe;
    assign coff[1950] = 64'h00005dd9ffffa8f4;
    assign coff[1951] = 64'h00005dd0ffffa8eb;
    assign coff[1952] = 64'h00005dc8ffffa8e2;
    assign coff[1953] = 64'h00005dbfffffa8d9;
    assign coff[1954] = 64'h00005db7ffffa8d0;
    assign coff[1955] = 64'h00005daeffffa8c6;
    assign coff[1956] = 64'h00005da5ffffa8bd;
    assign coff[1957] = 64'h00005d9dffffa8b4;
    assign coff[1958] = 64'h00005d94ffffa8ab;
    assign coff[1959] = 64'h00005d8cffffa8a2;
    assign coff[1960] = 64'h00005d83ffffa899;
    assign coff[1961] = 64'h00005d7affffa88f;
    assign coff[1962] = 64'h00005d72ffffa886;
    assign coff[1963] = 64'h00005d69ffffa87d;
    assign coff[1964] = 64'h00005d61ffffa874;
    assign coff[1965] = 64'h00005d58ffffa86b;
    assign coff[1966] = 64'h00005d50ffffa861;
    assign coff[1967] = 64'h00005d47ffffa858;
    assign coff[1968] = 64'h00005d3effffa84f;
    assign coff[1969] = 64'h00005d36ffffa846;
    assign coff[1970] = 64'h00005d2dffffa83d;
    assign coff[1971] = 64'h00005d24ffffa834;
    assign coff[1972] = 64'h00005d1cffffa82b;
    assign coff[1973] = 64'h00005d13ffffa821;
    assign coff[1974] = 64'h00005d0bffffa818;
    assign coff[1975] = 64'h00005d02ffffa80f;
    assign coff[1976] = 64'h00005cf9ffffa806;
    assign coff[1977] = 64'h00005cf1ffffa7fd;
    assign coff[1978] = 64'h00005ce8ffffa7f4;
    assign coff[1979] = 64'h00005cdfffffa7eb;
    assign coff[1980] = 64'h00005cd7ffffa7e2;
    assign coff[1981] = 64'h00005cceffffa7d8;
    assign coff[1982] = 64'h00005cc5ffffa7cf;
    assign coff[1983] = 64'h00005cbdffffa7c6;
    assign coff[1984] = 64'h00005cb4ffffa7bd;
    assign coff[1985] = 64'h00005cabffffa7b4;
    assign coff[1986] = 64'h00005ca3ffffa7ab;
    assign coff[1987] = 64'h00005c9affffa7a2;
    assign coff[1988] = 64'h00005c91ffffa799;
    assign coff[1989] = 64'h00005c89ffffa790;
    assign coff[1990] = 64'h00005c80ffffa787;
    assign coff[1991] = 64'h00005c77ffffa77e;
    assign coff[1992] = 64'h00005c6fffffa774;
    assign coff[1993] = 64'h00005c66ffffa76b;
    assign coff[1994] = 64'h00005c5dffffa762;
    assign coff[1995] = 64'h00005c55ffffa759;
    assign coff[1996] = 64'h00005c4cffffa750;
    assign coff[1997] = 64'h00005c43ffffa747;
    assign coff[1998] = 64'h00005c3affffa73e;
    assign coff[1999] = 64'h00005c32ffffa735;
    assign coff[2000] = 64'h00005c29ffffa72c;
    assign coff[2001] = 64'h00005c20ffffa723;
    assign coff[2002] = 64'h00005c18ffffa71a;
    assign coff[2003] = 64'h00005c0fffffa711;
    assign coff[2004] = 64'h00005c06ffffa708;
    assign coff[2005] = 64'h00005bfdffffa6ff;
    assign coff[2006] = 64'h00005bf5ffffa6f6;
    assign coff[2007] = 64'h00005becffffa6ed;
    assign coff[2008] = 64'h00005be3ffffa6e4;
    assign coff[2009] = 64'h00005bdaffffa6db;
    assign coff[2010] = 64'h00005bd2ffffa6d2;
    assign coff[2011] = 64'h00005bc9ffffa6c9;
    assign coff[2012] = 64'h00005bc0ffffa6c0;
    assign coff[2013] = 64'h00005bb7ffffa6b7;
    assign coff[2014] = 64'h00005bafffffa6ae;
    assign coff[2015] = 64'h00005ba6ffffa6a5;
    assign coff[2016] = 64'h00005b9dffffa69c;
    assign coff[2017] = 64'h00005b94ffffa693;
    assign coff[2018] = 64'h00005b8cffffa68a;
    assign coff[2019] = 64'h00005b83ffffa681;
    assign coff[2020] = 64'h00005b7affffa678;
    assign coff[2021] = 64'h00005b71ffffa66f;
    assign coff[2022] = 64'h00005b68ffffa666;
    assign coff[2023] = 64'h00005b60ffffa65d;
    assign coff[2024] = 64'h00005b57ffffa654;
    assign coff[2025] = 64'h00005b4effffa64b;
    assign coff[2026] = 64'h00005b45ffffa642;
    assign coff[2027] = 64'h00005b3cffffa639;
    assign coff[2028] = 64'h00005b34ffffa630;
    assign coff[2029] = 64'h00005b2bffffa627;
    assign coff[2030] = 64'h00005b22ffffa61e;
    assign coff[2031] = 64'h00005b19ffffa615;
    assign coff[2032] = 64'h00005b10ffffa60c;
    assign coff[2033] = 64'h00005b07ffffa603;
    assign coff[2034] = 64'h00005affffffa5fa;
    assign coff[2035] = 64'h00005af6ffffa5f1;
    assign coff[2036] = 64'h00005aedffffa5e8;
    assign coff[2037] = 64'h00005ae4ffffa5df;
    assign coff[2038] = 64'h00005adbffffa5d7;
    assign coff[2039] = 64'h00005ad2ffffa5ce;
    assign coff[2040] = 64'h00005ac9ffffa5c5;
    assign coff[2041] = 64'h00005ac1ffffa5bc;
    assign coff[2042] = 64'h00005ab8ffffa5b3;
    assign coff[2043] = 64'h00005aafffffa5aa;
    assign coff[2044] = 64'h00005aa6ffffa5a1;
    assign coff[2045] = 64'h00005a9dffffa598;
    assign coff[2046] = 64'h00005a94ffffa58f;
    assign coff[2047] = 64'h00005a8bffffa586;

    always_ff @(posedge clk, negedge rst_n) begin
        if(~rst_n) begin
            data_o_col1 <= 'b0;
            data_o_col2 <= 'b0;
        end else begin
            if ((addr_col1 == 'd0 || addr_col1 == 'd1024) && (valid == 1)) begin
                data_o_col1 <= coff[addr_col1];
                data_o_col2 <= 'b0;
            end else if(valid == 1) begin
                data_o_col1 <= coff[addr_col1];
                data_o_col2 <= coff[addr_col2];
            end else begin
                data_o_col1 <= 'b0;
                data_o_col2 <= 'b0;
            end       
        end
    end


endmodule