`timescale 1ns/1ps
module rom_2_rfft_data64
(
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic                     valid,
    input  logic [10:0]              addr_col1,
    input  logic [10:0]              addr_col2,
    output logic [63:0]              data_o_col1,
    output logic [63:0]              data_o_col2
);

    logic [63:0] coff[2047:0];

    assign coff[0   ] = 64'h00005a82ffffa57e;
    assign coff[1   ] = 64'h00005a7affffa575;
    assign coff[2   ] = 64'h00005a71ffffa56c;
    assign coff[3   ] = 64'h00005a68ffffa563;
    assign coff[4   ] = 64'h00005a5fffffa55a;
    assign coff[5   ] = 64'h00005a56ffffa551;
    assign coff[6   ] = 64'h00005a4dffffa548;
    assign coff[7   ] = 64'h00005a44ffffa53f;
    assign coff[8   ] = 64'h00005a3bffffa537;
    assign coff[9   ] = 64'h00005a32ffffa52e;
    assign coff[10  ] = 64'h00005a29ffffa525;
    assign coff[11  ] = 64'h00005a21ffffa51c;
    assign coff[12  ] = 64'h00005a18ffffa513;
    assign coff[13  ] = 64'h00005a0fffffa50a;
    assign coff[14  ] = 64'h00005a06ffffa501;
    assign coff[15  ] = 64'h000059fdffffa4f9;
    assign coff[16  ] = 64'h000059f4ffffa4f0;
    assign coff[17  ] = 64'h000059ebffffa4e7;
    assign coff[18  ] = 64'h000059e2ffffa4de;
    assign coff[19  ] = 64'h000059d9ffffa4d5;
    assign coff[20  ] = 64'h000059d0ffffa4cc;
    assign coff[21  ] = 64'h000059c7ffffa4c4;
    assign coff[22  ] = 64'h000059beffffa4bb;
    assign coff[23  ] = 64'h000059b5ffffa4b2;
    assign coff[24  ] = 64'h000059acffffa4a9;
    assign coff[25  ] = 64'h000059a3ffffa4a0;
    assign coff[26  ] = 64'h0000599affffa498;
    assign coff[27  ] = 64'h00005991ffffa48f;
    assign coff[28  ] = 64'h00005988ffffa486;
    assign coff[29  ] = 64'h0000597fffffa47d;
    assign coff[30  ] = 64'h00005976ffffa474;
    assign coff[31  ] = 64'h0000596dffffa46c;
    assign coff[32  ] = 64'h00005964ffffa463;
    assign coff[33  ] = 64'h0000595bffffa45a;
    assign coff[34  ] = 64'h00005952ffffa451;
    assign coff[35  ] = 64'h00005949ffffa449;
    assign coff[36  ] = 64'h00005940ffffa440;
    assign coff[37  ] = 64'h00005937ffffa437;
    assign coff[38  ] = 64'h0000592effffa42e;
    assign coff[39  ] = 64'h00005925ffffa426;
    assign coff[40  ] = 64'h0000591cffffa41d;
    assign coff[41  ] = 64'h00005913ffffa414;
    assign coff[42  ] = 64'h0000590affffa40b;
    assign coff[43  ] = 64'h00005901ffffa403;
    assign coff[44  ] = 64'h000058f8ffffa3fa;
    assign coff[45  ] = 64'h000058efffffa3f1;
    assign coff[46  ] = 64'h000058e6ffffa3e8;
    assign coff[47  ] = 64'h000058ddffffa3e0;
    assign coff[48  ] = 64'h000058d4ffffa3d7;
    assign coff[49  ] = 64'h000058cbffffa3ce;
    assign coff[50  ] = 64'h000058c2ffffa3c6;
    assign coff[51  ] = 64'h000058b9ffffa3bd;
    assign coff[52  ] = 64'h000058b0ffffa3b4;
    assign coff[53  ] = 64'h000058a7ffffa3ab;
    assign coff[54  ] = 64'h0000589effffa3a3;
    assign coff[55  ] = 64'h00005895ffffa39a;
    assign coff[56  ] = 64'h0000588cffffa391;
    assign coff[57  ] = 64'h00005882ffffa389;
    assign coff[58  ] = 64'h00005879ffffa380;
    assign coff[59  ] = 64'h00005870ffffa377;
    assign coff[60  ] = 64'h00005867ffffa36f;
    assign coff[61  ] = 64'h0000585effffa366;
    assign coff[62  ] = 64'h00005855ffffa35d;
    assign coff[63  ] = 64'h0000584cffffa355;
    assign coff[64  ] = 64'h00005843ffffa34c;
    assign coff[65  ] = 64'h0000583affffa343;
    assign coff[66  ] = 64'h00005831ffffa33b;
    assign coff[67  ] = 64'h00005828ffffa332;
    assign coff[68  ] = 64'h0000581effffa329;
    assign coff[69  ] = 64'h00005815ffffa321;
    assign coff[70  ] = 64'h0000580cffffa318;
    assign coff[71  ] = 64'h00005803ffffa30f;
    assign coff[72  ] = 64'h000057faffffa307;
    assign coff[73  ] = 64'h000057f1ffffa2fe;
    assign coff[74  ] = 64'h000057e8ffffa2f5;
    assign coff[75  ] = 64'h000057dfffffa2ed;
    assign coff[76  ] = 64'h000057d5ffffa2e4;
    assign coff[77  ] = 64'h000057ccffffa2dc;
    assign coff[78  ] = 64'h000057c3ffffa2d3;
    assign coff[79  ] = 64'h000057baffffa2ca;
    assign coff[80  ] = 64'h000057b1ffffa2c2;
    assign coff[81  ] = 64'h000057a8ffffa2b9;
    assign coff[82  ] = 64'h0000579fffffa2b0;
    assign coff[83  ] = 64'h00005795ffffa2a8;
    assign coff[84  ] = 64'h0000578cffffa29f;
    assign coff[85  ] = 64'h00005783ffffa297;
    assign coff[86  ] = 64'h0000577affffa28e;
    assign coff[87  ] = 64'h00005771ffffa286;
    assign coff[88  ] = 64'h00005767ffffa27d;
    assign coff[89  ] = 64'h0000575effffa274;
    assign coff[90  ] = 64'h00005755ffffa26c;
    assign coff[91  ] = 64'h0000574cffffa263;
    assign coff[92  ] = 64'h00005743ffffa25b;
    assign coff[93  ] = 64'h0000573affffa252;
    assign coff[94  ] = 64'h00005730ffffa249;
    assign coff[95  ] = 64'h00005727ffffa241;
    assign coff[96  ] = 64'h0000571effffa238;
    assign coff[97  ] = 64'h00005715ffffa230;
    assign coff[98  ] = 64'h0000570cffffa227;
    assign coff[99  ] = 64'h00005702ffffa21f;
    assign coff[100 ] = 64'h000056f9ffffa216;
    assign coff[101 ] = 64'h000056f0ffffa20e;
    assign coff[102 ] = 64'h000056e7ffffa205;
    assign coff[103 ] = 64'h000056ddffffa1fd;
    assign coff[104 ] = 64'h000056d4ffffa1f4;
    assign coff[105 ] = 64'h000056cbffffa1ec;
    assign coff[106 ] = 64'h000056c2ffffa1e3;
    assign coff[107 ] = 64'h000056b8ffffa1db;
    assign coff[108 ] = 64'h000056afffffa1d2;
    assign coff[109 ] = 64'h000056a6ffffa1c9;
    assign coff[110 ] = 64'h0000569dffffa1c1;
    assign coff[111 ] = 64'h00005693ffffa1b8;
    assign coff[112 ] = 64'h0000568affffa1b0;
    assign coff[113 ] = 64'h00005681ffffa1a8;
    assign coff[114 ] = 64'h00005678ffffa19f;
    assign coff[115 ] = 64'h0000566effffa197;
    assign coff[116 ] = 64'h00005665ffffa18e;
    assign coff[117 ] = 64'h0000565cffffa186;
    assign coff[118 ] = 64'h00005653ffffa17d;
    assign coff[119 ] = 64'h00005649ffffa175;
    assign coff[120 ] = 64'h00005640ffffa16c;
    assign coff[121 ] = 64'h00005637ffffa164;
    assign coff[122 ] = 64'h0000562dffffa15b;
    assign coff[123 ] = 64'h00005624ffffa153;
    assign coff[124 ] = 64'h0000561bffffa14a;
    assign coff[125 ] = 64'h00005612ffffa142;
    assign coff[126 ] = 64'h00005608ffffa139;
    assign coff[127 ] = 64'h000055ffffffa131;
    assign coff[128 ] = 64'h000055f6ffffa129;
    assign coff[129 ] = 64'h000055ecffffa120;
    assign coff[130 ] = 64'h000055e3ffffa118;
    assign coff[131 ] = 64'h000055daffffa10f;
    assign coff[132 ] = 64'h000055d0ffffa107;
    assign coff[133 ] = 64'h000055c7ffffa0fe;
    assign coff[134 ] = 64'h000055beffffa0f6;
    assign coff[135 ] = 64'h000055b4ffffa0ee;
    assign coff[136 ] = 64'h000055abffffa0e5;
    assign coff[137 ] = 64'h000055a2ffffa0dd;
    assign coff[138 ] = 64'h00005598ffffa0d4;
    assign coff[139 ] = 64'h0000558fffffa0cc;
    assign coff[140 ] = 64'h00005586ffffa0c4;
    assign coff[141 ] = 64'h0000557cffffa0bb;
    assign coff[142 ] = 64'h00005573ffffa0b3;
    assign coff[143 ] = 64'h0000556affffa0aa;
    assign coff[144 ] = 64'h00005560ffffa0a2;
    assign coff[145 ] = 64'h00005557ffffa09a;
    assign coff[146 ] = 64'h0000554effffa091;
    assign coff[147 ] = 64'h00005544ffffa089;
    assign coff[148 ] = 64'h0000553bffffa080;
    assign coff[149 ] = 64'h00005531ffffa078;
    assign coff[150 ] = 64'h00005528ffffa070;
    assign coff[151 ] = 64'h0000551fffffa067;
    assign coff[152 ] = 64'h00005515ffffa05f;
    assign coff[153 ] = 64'h0000550cffffa057;
    assign coff[154 ] = 64'h00005502ffffa04e;
    assign coff[155 ] = 64'h000054f9ffffa046;
    assign coff[156 ] = 64'h000054f0ffffa03e;
    assign coff[157 ] = 64'h000054e6ffffa035;
    assign coff[158 ] = 64'h000054ddffffa02d;
    assign coff[159 ] = 64'h000054d3ffffa025;
    assign coff[160 ] = 64'h000054caffffa01c;
    assign coff[161 ] = 64'h000054c1ffffa014;
    assign coff[162 ] = 64'h000054b7ffffa00c;
    assign coff[163 ] = 64'h000054aeffffa003;
    assign coff[164 ] = 64'h000054a4ffff9ffb;
    assign coff[165 ] = 64'h0000549bffff9ff3;
    assign coff[166 ] = 64'h00005491ffff9fea;
    assign coff[167 ] = 64'h00005488ffff9fe2;
    assign coff[168 ] = 64'h0000547fffff9fda;
    assign coff[169 ] = 64'h00005475ffff9fd2;
    assign coff[170 ] = 64'h0000546cffff9fc9;
    assign coff[171 ] = 64'h00005462ffff9fc1;
    assign coff[172 ] = 64'h00005459ffff9fb9;
    assign coff[173 ] = 64'h0000544fffff9fb0;
    assign coff[174 ] = 64'h00005446ffff9fa8;
    assign coff[175 ] = 64'h0000543cffff9fa0;
    assign coff[176 ] = 64'h00005433ffff9f98;
    assign coff[177 ] = 64'h0000542affff9f8f;
    assign coff[178 ] = 64'h00005420ffff9f87;
    assign coff[179 ] = 64'h00005417ffff9f7f;
    assign coff[180 ] = 64'h0000540dffff9f77;
    assign coff[181 ] = 64'h00005404ffff9f6e;
    assign coff[182 ] = 64'h000053faffff9f66;
    assign coff[183 ] = 64'h000053f1ffff9f5e;
    assign coff[184 ] = 64'h000053e7ffff9f56;
    assign coff[185 ] = 64'h000053deffff9f4d;
    assign coff[186 ] = 64'h000053d4ffff9f45;
    assign coff[187 ] = 64'h000053cbffff9f3d;
    assign coff[188 ] = 64'h000053c1ffff9f35;
    assign coff[189 ] = 64'h000053b8ffff9f2c;
    assign coff[190 ] = 64'h000053aeffff9f24;
    assign coff[191 ] = 64'h000053a5ffff9f1c;
    assign coff[192 ] = 64'h0000539bffff9f14;
    assign coff[193 ] = 64'h00005392ffff9f0c;
    assign coff[194 ] = 64'h00005388ffff9f03;
    assign coff[195 ] = 64'h0000537fffff9efb;
    assign coff[196 ] = 64'h00005375ffff9ef3;
    assign coff[197 ] = 64'h0000536cffff9eeb;
    assign coff[198 ] = 64'h00005362ffff9ee3;
    assign coff[199 ] = 64'h00005358ffff9eda;
    assign coff[200 ] = 64'h0000534fffff9ed2;
    assign coff[201 ] = 64'h00005345ffff9eca;
    assign coff[202 ] = 64'h0000533cffff9ec2;
    assign coff[203 ] = 64'h00005332ffff9eba;
    assign coff[204 ] = 64'h00005329ffff9eb2;
    assign coff[205 ] = 64'h0000531fffff9ea9;
    assign coff[206 ] = 64'h00005316ffff9ea1;
    assign coff[207 ] = 64'h0000530cffff9e99;
    assign coff[208 ] = 64'h00005303ffff9e91;
    assign coff[209 ] = 64'h000052f9ffff9e89;
    assign coff[210 ] = 64'h000052efffff9e81;
    assign coff[211 ] = 64'h000052e6ffff9e78;
    assign coff[212 ] = 64'h000052dcffff9e70;
    assign coff[213 ] = 64'h000052d3ffff9e68;
    assign coff[214 ] = 64'h000052c9ffff9e60;
    assign coff[215 ] = 64'h000052bfffff9e58;
    assign coff[216 ] = 64'h000052b6ffff9e50;
    assign coff[217 ] = 64'h000052acffff9e48;
    assign coff[218 ] = 64'h000052a3ffff9e40;
    assign coff[219 ] = 64'h00005299ffff9e37;
    assign coff[220 ] = 64'h00005290ffff9e2f;
    assign coff[221 ] = 64'h00005286ffff9e27;
    assign coff[222 ] = 64'h0000527cffff9e1f;
    assign coff[223 ] = 64'h00005273ffff9e17;
    assign coff[224 ] = 64'h00005269ffff9e0f;
    assign coff[225 ] = 64'h0000525fffff9e07;
    assign coff[226 ] = 64'h00005256ffff9dff;
    assign coff[227 ] = 64'h0000524cffff9df7;
    assign coff[228 ] = 64'h00005243ffff9def;
    assign coff[229 ] = 64'h00005239ffff9de7;
    assign coff[230 ] = 64'h0000522fffff9ddf;
    assign coff[231 ] = 64'h00005226ffff9dd6;
    assign coff[232 ] = 64'h0000521cffff9dce;
    assign coff[233 ] = 64'h00005212ffff9dc6;
    assign coff[234 ] = 64'h00005209ffff9dbe;
    assign coff[235 ] = 64'h000051ffffff9db6;
    assign coff[236 ] = 64'h000051f5ffff9dae;
    assign coff[237 ] = 64'h000051ecffff9da6;
    assign coff[238 ] = 64'h000051e2ffff9d9e;
    assign coff[239 ] = 64'h000051d8ffff9d96;
    assign coff[240 ] = 64'h000051cfffff9d8e;
    assign coff[241 ] = 64'h000051c5ffff9d86;
    assign coff[242 ] = 64'h000051bbffff9d7e;
    assign coff[243 ] = 64'h000051b2ffff9d76;
    assign coff[244 ] = 64'h000051a8ffff9d6e;
    assign coff[245 ] = 64'h0000519effff9d66;
    assign coff[246 ] = 64'h00005195ffff9d5e;
    assign coff[247 ] = 64'h0000518bffff9d56;
    assign coff[248 ] = 64'h00005181ffff9d4e;
    assign coff[249 ] = 64'h00005178ffff9d46;
    assign coff[250 ] = 64'h0000516effff9d3e;
    assign coff[251 ] = 64'h00005164ffff9d36;
    assign coff[252 ] = 64'h0000515bffff9d2e;
    assign coff[253 ] = 64'h00005151ffff9d26;
    assign coff[254 ] = 64'h00005147ffff9d1e;
    assign coff[255 ] = 64'h0000513effff9d16;
    assign coff[256 ] = 64'h00005134ffff9d0e;
    assign coff[257 ] = 64'h0000512affff9d06;
    assign coff[258 ] = 64'h00005120ffff9cfe;
    assign coff[259 ] = 64'h00005117ffff9cf6;
    assign coff[260 ] = 64'h0000510dffff9cee;
    assign coff[261 ] = 64'h00005103ffff9ce6;
    assign coff[262 ] = 64'h000050f9ffff9cde;
    assign coff[263 ] = 64'h000050f0ffff9cd6;
    assign coff[264 ] = 64'h000050e6ffff9cce;
    assign coff[265 ] = 64'h000050dcffff9cc6;
    assign coff[266 ] = 64'h000050d3ffff9cbe;
    assign coff[267 ] = 64'h000050c9ffff9cb7;
    assign coff[268 ] = 64'h000050bfffff9caf;
    assign coff[269 ] = 64'h000050b5ffff9ca7;
    assign coff[270 ] = 64'h000050acffff9c9f;
    assign coff[271 ] = 64'h000050a2ffff9c97;
    assign coff[272 ] = 64'h00005098ffff9c8f;
    assign coff[273 ] = 64'h0000508effff9c87;
    assign coff[274 ] = 64'h00005084ffff9c7f;
    assign coff[275 ] = 64'h0000507bffff9c77;
    assign coff[276 ] = 64'h00005071ffff9c6f;
    assign coff[277 ] = 64'h00005067ffff9c67;
    assign coff[278 ] = 64'h0000505dffff9c60;
    assign coff[279 ] = 64'h00005054ffff9c58;
    assign coff[280 ] = 64'h0000504affff9c50;
    assign coff[281 ] = 64'h00005040ffff9c48;
    assign coff[282 ] = 64'h00005036ffff9c40;
    assign coff[283 ] = 64'h0000502cffff9c38;
    assign coff[284 ] = 64'h00005023ffff9c30;
    assign coff[285 ] = 64'h00005019ffff9c28;
    assign coff[286 ] = 64'h0000500fffff9c21;
    assign coff[287 ] = 64'h00005005ffff9c19;
    assign coff[288 ] = 64'h00004ffbffff9c11;
    assign coff[289 ] = 64'h00004ff2ffff9c09;
    assign coff[290 ] = 64'h00004fe8ffff9c01;
    assign coff[291 ] = 64'h00004fdeffff9bf9;
    assign coff[292 ] = 64'h00004fd4ffff9bf1;
    assign coff[293 ] = 64'h00004fcaffff9bea;
    assign coff[294 ] = 64'h00004fc0ffff9be2;
    assign coff[295 ] = 64'h00004fb7ffff9bda;
    assign coff[296 ] = 64'h00004fadffff9bd2;
    assign coff[297 ] = 64'h00004fa3ffff9bca;
    assign coff[298 ] = 64'h00004f99ffff9bc2;
    assign coff[299 ] = 64'h00004f8fffff9bbb;
    assign coff[300 ] = 64'h00004f85ffff9bb3;
    assign coff[301 ] = 64'h00004f7cffff9bab;
    assign coff[302 ] = 64'h00004f72ffff9ba3;
    assign coff[303 ] = 64'h00004f68ffff9b9b;
    assign coff[304 ] = 64'h00004f5effff9b94;
    assign coff[305 ] = 64'h00004f54ffff9b8c;
    assign coff[306 ] = 64'h00004f4affff9b84;
    assign coff[307 ] = 64'h00004f40ffff9b7c;
    assign coff[308 ] = 64'h00004f37ffff9b75;
    assign coff[309 ] = 64'h00004f2dffff9b6d;
    assign coff[310 ] = 64'h00004f23ffff9b65;
    assign coff[311 ] = 64'h00004f19ffff9b5d;
    assign coff[312 ] = 64'h00004f0fffff9b55;
    assign coff[313 ] = 64'h00004f05ffff9b4e;
    assign coff[314 ] = 64'h00004efbffff9b46;
    assign coff[315 ] = 64'h00004ef1ffff9b3e;
    assign coff[316 ] = 64'h00004ee8ffff9b36;
    assign coff[317 ] = 64'h00004edeffff9b2f;
    assign coff[318 ] = 64'h00004ed4ffff9b27;
    assign coff[319 ] = 64'h00004ecaffff9b1f;
    assign coff[320 ] = 64'h00004ec0ffff9b17;
    assign coff[321 ] = 64'h00004eb6ffff9b10;
    assign coff[322 ] = 64'h00004eacffff9b08;
    assign coff[323 ] = 64'h00004ea2ffff9b00;
    assign coff[324 ] = 64'h00004e98ffff9af9;
    assign coff[325 ] = 64'h00004e8effff9af1;
    assign coff[326 ] = 64'h00004e84ffff9ae9;
    assign coff[327 ] = 64'h00004e7affff9ae1;
    assign coff[328 ] = 64'h00004e71ffff9ada;
    assign coff[329 ] = 64'h00004e67ffff9ad2;
    assign coff[330 ] = 64'h00004e5dffff9aca;
    assign coff[331 ] = 64'h00004e53ffff9ac3;
    assign coff[332 ] = 64'h00004e49ffff9abb;
    assign coff[333 ] = 64'h00004e3fffff9ab3;
    assign coff[334 ] = 64'h00004e35ffff9aac;
    assign coff[335 ] = 64'h00004e2bffff9aa4;
    assign coff[336 ] = 64'h00004e21ffff9a9c;
    assign coff[337 ] = 64'h00004e17ffff9a95;
    assign coff[338 ] = 64'h00004e0dffff9a8d;
    assign coff[339 ] = 64'h00004e03ffff9a85;
    assign coff[340 ] = 64'h00004df9ffff9a7e;
    assign coff[341 ] = 64'h00004defffff9a76;
    assign coff[342 ] = 64'h00004de5ffff9a6e;
    assign coff[343 ] = 64'h00004ddbffff9a67;
    assign coff[344 ] = 64'h00004dd1ffff9a5f;
    assign coff[345 ] = 64'h00004dc7ffff9a57;
    assign coff[346 ] = 64'h00004dbdffff9a50;
    assign coff[347 ] = 64'h00004db3ffff9a48;
    assign coff[348 ] = 64'h00004da9ffff9a40;
    assign coff[349 ] = 64'h00004d9fffff9a39;
    assign coff[350 ] = 64'h00004d95ffff9a31;
    assign coff[351 ] = 64'h00004d8bffff9a2a;
    assign coff[352 ] = 64'h00004d81ffff9a22;
    assign coff[353 ] = 64'h00004d77ffff9a1a;
    assign coff[354 ] = 64'h00004d6dffff9a13;
    assign coff[355 ] = 64'h00004d63ffff9a0b;
    assign coff[356 ] = 64'h00004d59ffff9a04;
    assign coff[357 ] = 64'h00004d4fffff99fc;
    assign coff[358 ] = 64'h00004d45ffff99f4;
    assign coff[359 ] = 64'h00004d3bffff99ed;
    assign coff[360 ] = 64'h00004d31ffff99e5;
    assign coff[361 ] = 64'h00004d27ffff99de;
    assign coff[362 ] = 64'h00004d1dffff99d6;
    assign coff[363 ] = 64'h00004d13ffff99cf;
    assign coff[364 ] = 64'h00004d09ffff99c7;
    assign coff[365 ] = 64'h00004cffffff99bf;
    assign coff[366 ] = 64'h00004cf5ffff99b8;
    assign coff[367 ] = 64'h00004cebffff99b0;
    assign coff[368 ] = 64'h00004ce1ffff99a9;
    assign coff[369 ] = 64'h00004cd7ffff99a1;
    assign coff[370 ] = 64'h00004ccdffff999a;
    assign coff[371 ] = 64'h00004cc3ffff9992;
    assign coff[372 ] = 64'h00004cb9ffff998b;
    assign coff[373 ] = 64'h00004cafffff9983;
    assign coff[374 ] = 64'h00004ca5ffff997c;
    assign coff[375 ] = 64'h00004c9bffff9974;
    assign coff[376 ] = 64'h00004c91ffff996d;
    assign coff[377 ] = 64'h00004c86ffff9965;
    assign coff[378 ] = 64'h00004c7cffff995d;
    assign coff[379 ] = 64'h00004c72ffff9956;
    assign coff[380 ] = 64'h00004c68ffff994e;
    assign coff[381 ] = 64'h00004c5effff9947;
    assign coff[382 ] = 64'h00004c54ffff993f;
    assign coff[383 ] = 64'h00004c4affff9938;
    assign coff[384 ] = 64'h00004c40ffff9930;
    assign coff[385 ] = 64'h00004c36ffff9929;
    assign coff[386 ] = 64'h00004c2cffff9922;
    assign coff[387 ] = 64'h00004c22ffff991a;
    assign coff[388 ] = 64'h00004c17ffff9913;
    assign coff[389 ] = 64'h00004c0dffff990b;
    assign coff[390 ] = 64'h00004c03ffff9904;
    assign coff[391 ] = 64'h00004bf9ffff98fc;
    assign coff[392 ] = 64'h00004befffff98f5;
    assign coff[393 ] = 64'h00004be5ffff98ed;
    assign coff[394 ] = 64'h00004bdbffff98e6;
    assign coff[395 ] = 64'h00004bd1ffff98de;
    assign coff[396 ] = 64'h00004bc7ffff98d7;
    assign coff[397 ] = 64'h00004bbcffff98d0;
    assign coff[398 ] = 64'h00004bb2ffff98c8;
    assign coff[399 ] = 64'h00004ba8ffff98c1;
    assign coff[400 ] = 64'h00004b9effff98b9;
    assign coff[401 ] = 64'h00004b94ffff98b2;
    assign coff[402 ] = 64'h00004b8affff98aa;
    assign coff[403 ] = 64'h00004b80ffff98a3;
    assign coff[404 ] = 64'h00004b75ffff989c;
    assign coff[405 ] = 64'h00004b6bffff9894;
    assign coff[406 ] = 64'h00004b61ffff988d;
    assign coff[407 ] = 64'h00004b57ffff9885;
    assign coff[408 ] = 64'h00004b4dffff987e;
    assign coff[409 ] = 64'h00004b43ffff9877;
    assign coff[410 ] = 64'h00004b38ffff986f;
    assign coff[411 ] = 64'h00004b2effff9868;
    assign coff[412 ] = 64'h00004b24ffff9860;
    assign coff[413 ] = 64'h00004b1affff9859;
    assign coff[414 ] = 64'h00004b10ffff9852;
    assign coff[415 ] = 64'h00004b06ffff984a;
    assign coff[416 ] = 64'h00004afbffff9843;
    assign coff[417 ] = 64'h00004af1ffff983c;
    assign coff[418 ] = 64'h00004ae7ffff9834;
    assign coff[419 ] = 64'h00004addffff982d;
    assign coff[420 ] = 64'h00004ad3ffff9826;
    assign coff[421 ] = 64'h00004ac8ffff981e;
    assign coff[422 ] = 64'h00004abeffff9817;
    assign coff[423 ] = 64'h00004ab4ffff9810;
    assign coff[424 ] = 64'h00004aaaffff9808;
    assign coff[425 ] = 64'h00004aa0ffff9801;
    assign coff[426 ] = 64'h00004a95ffff97fa;
    assign coff[427 ] = 64'h00004a8bffff97f2;
    assign coff[428 ] = 64'h00004a81ffff97eb;
    assign coff[429 ] = 64'h00004a77ffff97e4;
    assign coff[430 ] = 64'h00004a6dffff97dc;
    assign coff[431 ] = 64'h00004a62ffff97d5;
    assign coff[432 ] = 64'h00004a58ffff97ce;
    assign coff[433 ] = 64'h00004a4effff97c6;
    assign coff[434 ] = 64'h00004a44ffff97bf;
    assign coff[435 ] = 64'h00004a39ffff97b8;
    assign coff[436 ] = 64'h00004a2fffff97b0;
    assign coff[437 ] = 64'h00004a25ffff97a9;
    assign coff[438 ] = 64'h00004a1bffff97a2;
    assign coff[439 ] = 64'h00004a10ffff979b;
    assign coff[440 ] = 64'h00004a06ffff9793;
    assign coff[441 ] = 64'h000049fcffff978c;
    assign coff[442 ] = 64'h000049f2ffff9785;
    assign coff[443 ] = 64'h000049e7ffff977e;
    assign coff[444 ] = 64'h000049ddffff9776;
    assign coff[445 ] = 64'h000049d3ffff976f;
    assign coff[446 ] = 64'h000049c9ffff9768;
    assign coff[447 ] = 64'h000049beffff9761;
    assign coff[448 ] = 64'h000049b4ffff9759;
    assign coff[449 ] = 64'h000049aaffff9752;
    assign coff[450 ] = 64'h000049a0ffff974b;
    assign coff[451 ] = 64'h00004995ffff9744;
    assign coff[452 ] = 64'h0000498bffff973c;
    assign coff[453 ] = 64'h00004981ffff9735;
    assign coff[454 ] = 64'h00004976ffff972e;
    assign coff[455 ] = 64'h0000496cffff9727;
    assign coff[456 ] = 64'h00004962ffff9720;
    assign coff[457 ] = 64'h00004958ffff9718;
    assign coff[458 ] = 64'h0000494dffff9711;
    assign coff[459 ] = 64'h00004943ffff970a;
    assign coff[460 ] = 64'h00004939ffff9703;
    assign coff[461 ] = 64'h0000492effff96fc;
    assign coff[462 ] = 64'h00004924ffff96f4;
    assign coff[463 ] = 64'h0000491affff96ed;
    assign coff[464 ] = 64'h0000490fffff96e6;
    assign coff[465 ] = 64'h00004905ffff96df;
    assign coff[466 ] = 64'h000048fbffff96d8;
    assign coff[467 ] = 64'h000048f0ffff96d1;
    assign coff[468 ] = 64'h000048e6ffff96c9;
    assign coff[469 ] = 64'h000048dcffff96c2;
    assign coff[470 ] = 64'h000048d1ffff96bb;
    assign coff[471 ] = 64'h000048c7ffff96b4;
    assign coff[472 ] = 64'h000048bdffff96ad;
    assign coff[473 ] = 64'h000048b2ffff96a6;
    assign coff[474 ] = 64'h000048a8ffff969f;
    assign coff[475 ] = 64'h0000489effff9697;
    assign coff[476 ] = 64'h00004893ffff9690;
    assign coff[477 ] = 64'h00004889ffff9689;
    assign coff[478 ] = 64'h0000487fffff9682;
    assign coff[479 ] = 64'h00004874ffff967b;
    assign coff[480 ] = 64'h0000486affff9674;
    assign coff[481 ] = 64'h00004860ffff966d;
    assign coff[482 ] = 64'h00004855ffff9666;
    assign coff[483 ] = 64'h0000484bffff965f;
    assign coff[484 ] = 64'h00004840ffff9657;
    assign coff[485 ] = 64'h00004836ffff9650;
    assign coff[486 ] = 64'h0000482cffff9649;
    assign coff[487 ] = 64'h00004821ffff9642;
    assign coff[488 ] = 64'h00004817ffff963b;
    assign coff[489 ] = 64'h0000480dffff9634;
    assign coff[490 ] = 64'h00004802ffff962d;
    assign coff[491 ] = 64'h000047f8ffff9626;
    assign coff[492 ] = 64'h000047edffff961f;
    assign coff[493 ] = 64'h000047e3ffff9618;
    assign coff[494 ] = 64'h000047d9ffff9611;
    assign coff[495 ] = 64'h000047ceffff960a;
    assign coff[496 ] = 64'h000047c4ffff9603;
    assign coff[497 ] = 64'h000047b9ffff95fc;
    assign coff[498 ] = 64'h000047afffff95f5;
    assign coff[499 ] = 64'h000047a5ffff95ee;
    assign coff[500 ] = 64'h0000479affff95e6;
    assign coff[501 ] = 64'h00004790ffff95df;
    assign coff[502 ] = 64'h00004785ffff95d8;
    assign coff[503 ] = 64'h0000477bffff95d1;
    assign coff[504 ] = 64'h00004770ffff95ca;
    assign coff[505 ] = 64'h00004766ffff95c3;
    assign coff[506 ] = 64'h0000475cffff95bc;
    assign coff[507 ] = 64'h00004751ffff95b5;
    assign coff[508 ] = 64'h00004747ffff95ae;
    assign coff[509 ] = 64'h0000473cffff95a7;
    assign coff[510 ] = 64'h00004732ffff95a0;
    assign coff[511 ] = 64'h00004727ffff9599;
    assign coff[512 ] = 64'h0000471dffff9592;
    assign coff[513 ] = 64'h00004712ffff958b;
    assign coff[514 ] = 64'h00004708ffff9584;
    assign coff[515 ] = 64'h000046feffff957d;
    assign coff[516 ] = 64'h000046f3ffff9577;
    assign coff[517 ] = 64'h000046e9ffff9570;
    assign coff[518 ] = 64'h000046deffff9569;
    assign coff[519 ] = 64'h000046d4ffff9562;
    assign coff[520 ] = 64'h000046c9ffff955b;
    assign coff[521 ] = 64'h000046bfffff9554;
    assign coff[522 ] = 64'h000046b4ffff954d;
    assign coff[523 ] = 64'h000046aaffff9546;
    assign coff[524 ] = 64'h0000469fffff953f;
    assign coff[525 ] = 64'h00004695ffff9538;
    assign coff[526 ] = 64'h0000468affff9531;
    assign coff[527 ] = 64'h00004680ffff952a;
    assign coff[528 ] = 64'h00004675ffff9523;
    assign coff[529 ] = 64'h0000466bffff951c;
    assign coff[530 ] = 64'h00004660ffff9515;
    assign coff[531 ] = 64'h00004656ffff950e;
    assign coff[532 ] = 64'h0000464bffff9508;
    assign coff[533 ] = 64'h00004641ffff9501;
    assign coff[534 ] = 64'h00004636ffff94fa;
    assign coff[535 ] = 64'h0000462cffff94f3;
    assign coff[536 ] = 64'h00004621ffff94ec;
    assign coff[537 ] = 64'h00004617ffff94e5;
    assign coff[538 ] = 64'h0000460cffff94de;
    assign coff[539 ] = 64'h00004602ffff94d7;
    assign coff[540 ] = 64'h000045f7ffff94d0;
    assign coff[541 ] = 64'h000045edffff94ca;
    assign coff[542 ] = 64'h000045e2ffff94c3;
    assign coff[543 ] = 64'h000045d8ffff94bc;
    assign coff[544 ] = 64'h000045cdffff94b5;
    assign coff[545 ] = 64'h000045c3ffff94ae;
    assign coff[546 ] = 64'h000045b8ffff94a7;
    assign coff[547 ] = 64'h000045aeffff94a1;
    assign coff[548 ] = 64'h000045a3ffff949a;
    assign coff[549 ] = 64'h00004599ffff9493;
    assign coff[550 ] = 64'h0000458effff948c;
    assign coff[551 ] = 64'h00004583ffff9485;
    assign coff[552 ] = 64'h00004579ffff947e;
    assign coff[553 ] = 64'h0000456effff9478;
    assign coff[554 ] = 64'h00004564ffff9471;
    assign coff[555 ] = 64'h00004559ffff946a;
    assign coff[556 ] = 64'h0000454fffff9463;
    assign coff[557 ] = 64'h00004544ffff945c;
    assign coff[558 ] = 64'h00004539ffff9456;
    assign coff[559 ] = 64'h0000452fffff944f;
    assign coff[560 ] = 64'h00004524ffff9448;
    assign coff[561 ] = 64'h0000451affff9441;
    assign coff[562 ] = 64'h0000450fffff943a;
    assign coff[563 ] = 64'h00004505ffff9434;
    assign coff[564 ] = 64'h000044faffff942d;
    assign coff[565 ] = 64'h000044efffff9426;
    assign coff[566 ] = 64'h000044e5ffff941f;
    assign coff[567 ] = 64'h000044daffff9419;
    assign coff[568 ] = 64'h000044d0ffff9412;
    assign coff[569 ] = 64'h000044c5ffff940b;
    assign coff[570 ] = 64'h000044baffff9404;
    assign coff[571 ] = 64'h000044b0ffff93fe;
    assign coff[572 ] = 64'h000044a5ffff93f7;
    assign coff[573 ] = 64'h0000449bffff93f0;
    assign coff[574 ] = 64'h00004490ffff93e9;
    assign coff[575 ] = 64'h00004485ffff93e3;
    assign coff[576 ] = 64'h0000447bffff93dc;
    assign coff[577 ] = 64'h00004470ffff93d5;
    assign coff[578 ] = 64'h00004466ffff93ce;
    assign coff[579 ] = 64'h0000445bffff93c8;
    assign coff[580 ] = 64'h00004450ffff93c1;
    assign coff[581 ] = 64'h00004446ffff93ba;
    assign coff[582 ] = 64'h0000443bffff93b4;
    assign coff[583 ] = 64'h00004430ffff93ad;
    assign coff[584 ] = 64'h00004426ffff93a6;
    assign coff[585 ] = 64'h0000441bffff939f;
    assign coff[586 ] = 64'h00004411ffff9399;
    assign coff[587 ] = 64'h00004406ffff9392;
    assign coff[588 ] = 64'h000043fbffff938b;
    assign coff[589 ] = 64'h000043f1ffff9385;
    assign coff[590 ] = 64'h000043e6ffff937e;
    assign coff[591 ] = 64'h000043dbffff9377;
    assign coff[592 ] = 64'h000043d1ffff9371;
    assign coff[593 ] = 64'h000043c6ffff936a;
    assign coff[594 ] = 64'h000043bbffff9363;
    assign coff[595 ] = 64'h000043b1ffff935d;
    assign coff[596 ] = 64'h000043a6ffff9356;
    assign coff[597 ] = 64'h0000439bffff9350;
    assign coff[598 ] = 64'h00004391ffff9349;
    assign coff[599 ] = 64'h00004386ffff9342;
    assign coff[600 ] = 64'h0000437bffff933c;
    assign coff[601 ] = 64'h00004371ffff9335;
    assign coff[602 ] = 64'h00004366ffff932e;
    assign coff[603 ] = 64'h0000435bffff9328;
    assign coff[604 ] = 64'h00004351ffff9321;
    assign coff[605 ] = 64'h00004346ffff931b;
    assign coff[606 ] = 64'h0000433bffff9314;
    assign coff[607 ] = 64'h00004330ffff930d;
    assign coff[608 ] = 64'h00004326ffff9307;
    assign coff[609 ] = 64'h0000431bffff9300;
    assign coff[610 ] = 64'h00004310ffff92fa;
    assign coff[611 ] = 64'h00004306ffff92f3;
    assign coff[612 ] = 64'h000042fbffff92ec;
    assign coff[613 ] = 64'h000042f0ffff92e6;
    assign coff[614 ] = 64'h000042e6ffff92df;
    assign coff[615 ] = 64'h000042dbffff92d9;
    assign coff[616 ] = 64'h000042d0ffff92d2;
    assign coff[617 ] = 64'h000042c5ffff92cc;
    assign coff[618 ] = 64'h000042bbffff92c5;
    assign coff[619 ] = 64'h000042b0ffff92bf;
    assign coff[620 ] = 64'h000042a5ffff92b8;
    assign coff[621 ] = 64'h0000429affff92b1;
    assign coff[622 ] = 64'h00004290ffff92ab;
    assign coff[623 ] = 64'h00004285ffff92a4;
    assign coff[624 ] = 64'h0000427affff929e;
    assign coff[625 ] = 64'h00004270ffff9297;
    assign coff[626 ] = 64'h00004265ffff9291;
    assign coff[627 ] = 64'h0000425affff928a;
    assign coff[628 ] = 64'h0000424fffff9284;
    assign coff[629 ] = 64'h00004245ffff927d;
    assign coff[630 ] = 64'h0000423affff9277;
    assign coff[631 ] = 64'h0000422fffff9270;
    assign coff[632 ] = 64'h00004224ffff926a;
    assign coff[633 ] = 64'h0000421affff9263;
    assign coff[634 ] = 64'h0000420fffff925d;
    assign coff[635 ] = 64'h00004204ffff9256;
    assign coff[636 ] = 64'h000041f9ffff9250;
    assign coff[637 ] = 64'h000041eeffff9249;
    assign coff[638 ] = 64'h000041e4ffff9243;
    assign coff[639 ] = 64'h000041d9ffff923c;
    assign coff[640 ] = 64'h000041ceffff9236;
    assign coff[641 ] = 64'h000041c3ffff922f;
    assign coff[642 ] = 64'h000041b9ffff9229;
    assign coff[643 ] = 64'h000041aeffff9223;
    assign coff[644 ] = 64'h000041a3ffff921c;
    assign coff[645 ] = 64'h00004198ffff9216;
    assign coff[646 ] = 64'h0000418dffff920f;
    assign coff[647 ] = 64'h00004183ffff9209;
    assign coff[648 ] = 64'h00004178ffff9202;
    assign coff[649 ] = 64'h0000416dffff91fc;
    assign coff[650 ] = 64'h00004162ffff91f6;
    assign coff[651 ] = 64'h00004157ffff91ef;
    assign coff[652 ] = 64'h0000414dffff91e9;
    assign coff[653 ] = 64'h00004142ffff91e2;
    assign coff[654 ] = 64'h00004137ffff91dc;
    assign coff[655 ] = 64'h0000412cffff91d6;
    assign coff[656 ] = 64'h00004121ffff91cf;
    assign coff[657 ] = 64'h00004117ffff91c9;
    assign coff[658 ] = 64'h0000410cffff91c2;
    assign coff[659 ] = 64'h00004101ffff91bc;
    assign coff[660 ] = 64'h000040f6ffff91b6;
    assign coff[661 ] = 64'h000040ebffff91af;
    assign coff[662 ] = 64'h000040e0ffff91a9;
    assign coff[663 ] = 64'h000040d6ffff91a2;
    assign coff[664 ] = 64'h000040cbffff919c;
    assign coff[665 ] = 64'h000040c0ffff9196;
    assign coff[666 ] = 64'h000040b5ffff918f;
    assign coff[667 ] = 64'h000040aaffff9189;
    assign coff[668 ] = 64'h0000409fffff9183;
    assign coff[669 ] = 64'h00004095ffff917c;
    assign coff[670 ] = 64'h0000408affff9176;
    assign coff[671 ] = 64'h0000407fffff9170;
    assign coff[672 ] = 64'h00004074ffff9169;
    assign coff[673 ] = 64'h00004069ffff9163;
    assign coff[674 ] = 64'h0000405effff915d;
    assign coff[675 ] = 64'h00004053ffff9156;
    assign coff[676 ] = 64'h00004048ffff9150;
    assign coff[677 ] = 64'h0000403effff914a;
    assign coff[678 ] = 64'h00004033ffff9143;
    assign coff[679 ] = 64'h00004028ffff913d;
    assign coff[680 ] = 64'h0000401dffff9137;
    assign coff[681 ] = 64'h00004012ffff9131;
    assign coff[682 ] = 64'h00004007ffff912a;
    assign coff[683 ] = 64'h00003ffcffff9124;
    assign coff[684 ] = 64'h00003ff1ffff911e;
    assign coff[685 ] = 64'h00003fe7ffff9117;
    assign coff[686 ] = 64'h00003fdcffff9111;
    assign coff[687 ] = 64'h00003fd1ffff910b;
    assign coff[688 ] = 64'h00003fc6ffff9105;
    assign coff[689 ] = 64'h00003fbbffff90fe;
    assign coff[690 ] = 64'h00003fb0ffff90f8;
    assign coff[691 ] = 64'h00003fa5ffff90f2;
    assign coff[692 ] = 64'h00003f9affff90ec;
    assign coff[693 ] = 64'h00003f8fffff90e5;
    assign coff[694 ] = 64'h00003f85ffff90df;
    assign coff[695 ] = 64'h00003f7affff90d9;
    assign coff[696 ] = 64'h00003f6fffff90d3;
    assign coff[697 ] = 64'h00003f64ffff90cc;
    assign coff[698 ] = 64'h00003f59ffff90c6;
    assign coff[699 ] = 64'h00003f4effff90c0;
    assign coff[700 ] = 64'h00003f43ffff90ba;
    assign coff[701 ] = 64'h00003f38ffff90b4;
    assign coff[702 ] = 64'h00003f2dffff90ad;
    assign coff[703 ] = 64'h00003f22ffff90a7;
    assign coff[704 ] = 64'h00003f17ffff90a1;
    assign coff[705 ] = 64'h00003f0cffff909b;
    assign coff[706 ] = 64'h00003f01ffff9095;
    assign coff[707 ] = 64'h00003ef6ffff908e;
    assign coff[708 ] = 64'h00003eecffff9088;
    assign coff[709 ] = 64'h00003ee1ffff9082;
    assign coff[710 ] = 64'h00003ed6ffff907c;
    assign coff[711 ] = 64'h00003ecbffff9076;
    assign coff[712 ] = 64'h00003ec0ffff9070;
    assign coff[713 ] = 64'h00003eb5ffff9069;
    assign coff[714 ] = 64'h00003eaaffff9063;
    assign coff[715 ] = 64'h00003e9fffff905d;
    assign coff[716 ] = 64'h00003e94ffff9057;
    assign coff[717 ] = 64'h00003e89ffff9051;
    assign coff[718 ] = 64'h00003e7effff904b;
    assign coff[719 ] = 64'h00003e73ffff9045;
    assign coff[720 ] = 64'h00003e68ffff903e;
    assign coff[721 ] = 64'h00003e5dffff9038;
    assign coff[722 ] = 64'h00003e52ffff9032;
    assign coff[723 ] = 64'h00003e47ffff902c;
    assign coff[724 ] = 64'h00003e3cffff9026;
    assign coff[725 ] = 64'h00003e31ffff9020;
    assign coff[726 ] = 64'h00003e26ffff901a;
    assign coff[727 ] = 64'h00003e1bffff9014;
    assign coff[728 ] = 64'h00003e10ffff900e;
    assign coff[729 ] = 64'h00003e05ffff9007;
    assign coff[730 ] = 64'h00003dfaffff9001;
    assign coff[731 ] = 64'h00003defffff8ffb;
    assign coff[732 ] = 64'h00003de4ffff8ff5;
    assign coff[733 ] = 64'h00003dd9ffff8fef;
    assign coff[734 ] = 64'h00003dceffff8fe9;
    assign coff[735 ] = 64'h00003dc3ffff8fe3;
    assign coff[736 ] = 64'h00003db8ffff8fdd;
    assign coff[737 ] = 64'h00003dadffff8fd7;
    assign coff[738 ] = 64'h00003da2ffff8fd1;
    assign coff[739 ] = 64'h00003d97ffff8fcb;
    assign coff[740 ] = 64'h00003d8cffff8fc5;
    assign coff[741 ] = 64'h00003d81ffff8fbf;
    assign coff[742 ] = 64'h00003d76ffff8fb9;
    assign coff[743 ] = 64'h00003d6bffff8fb3;
    assign coff[744 ] = 64'h00003d60ffff8fad;
    assign coff[745 ] = 64'h00003d55ffff8fa7;
    assign coff[746 ] = 64'h00003d4affff8fa1;
    assign coff[747 ] = 64'h00003d3fffff8f9b;
    assign coff[748 ] = 64'h00003d34ffff8f95;
    assign coff[749 ] = 64'h00003d29ffff8f8f;
    assign coff[750 ] = 64'h00003d1effff8f89;
    assign coff[751 ] = 64'h00003d13ffff8f83;
    assign coff[752 ] = 64'h00003d08ffff8f7d;
    assign coff[753 ] = 64'h00003cfdffff8f77;
    assign coff[754 ] = 64'h00003cf2ffff8f71;
    assign coff[755 ] = 64'h00003ce7ffff8f6b;
    assign coff[756 ] = 64'h00003cdcffff8f65;
    assign coff[757 ] = 64'h00003cd0ffff8f5f;
    assign coff[758 ] = 64'h00003cc5ffff8f59;
    assign coff[759 ] = 64'h00003cbaffff8f53;
    assign coff[760 ] = 64'h00003cafffff8f4d;
    assign coff[761 ] = 64'h00003ca4ffff8f47;
    assign coff[762 ] = 64'h00003c99ffff8f41;
    assign coff[763 ] = 64'h00003c8effff8f3b;
    assign coff[764 ] = 64'h00003c83ffff8f35;
    assign coff[765 ] = 64'h00003c78ffff8f2f;
    assign coff[766 ] = 64'h00003c6dffff8f29;
    assign coff[767 ] = 64'h00003c62ffff8f23;
    assign coff[768 ] = 64'h00003c57ffff8f1d;
    assign coff[769 ] = 64'h00003c4cffff8f17;
    assign coff[770 ] = 64'h00003c41ffff8f11;
    assign coff[771 ] = 64'h00003c35ffff8f0b;
    assign coff[772 ] = 64'h00003c2affff8f06;
    assign coff[773 ] = 64'h00003c1fffff8f00;
    assign coff[774 ] = 64'h00003c14ffff8efa;
    assign coff[775 ] = 64'h00003c09ffff8ef4;
    assign coff[776 ] = 64'h00003bfeffff8eee;
    assign coff[777 ] = 64'h00003bf3ffff8ee8;
    assign coff[778 ] = 64'h00003be8ffff8ee2;
    assign coff[779 ] = 64'h00003bddffff8edc;
    assign coff[780 ] = 64'h00003bd2ffff8ed6;
    assign coff[781 ] = 64'h00003bc6ffff8ed1;
    assign coff[782 ] = 64'h00003bbbffff8ecb;
    assign coff[783 ] = 64'h00003bb0ffff8ec5;
    assign coff[784 ] = 64'h00003ba5ffff8ebf;
    assign coff[785 ] = 64'h00003b9affff8eb9;
    assign coff[786 ] = 64'h00003b8fffff8eb3;
    assign coff[787 ] = 64'h00003b84ffff8ead;
    assign coff[788 ] = 64'h00003b79ffff8ea8;
    assign coff[789 ] = 64'h00003b6dffff8ea2;
    assign coff[790 ] = 64'h00003b62ffff8e9c;
    assign coff[791 ] = 64'h00003b57ffff8e96;
    assign coff[792 ] = 64'h00003b4cffff8e90;
    assign coff[793 ] = 64'h00003b41ffff8e8a;
    assign coff[794 ] = 64'h00003b36ffff8e85;
    assign coff[795 ] = 64'h00003b2bffff8e7f;
    assign coff[796 ] = 64'h00003b20ffff8e79;
    assign coff[797 ] = 64'h00003b14ffff8e73;
    assign coff[798 ] = 64'h00003b09ffff8e6d;
    assign coff[799 ] = 64'h00003afeffff8e68;
    assign coff[800 ] = 64'h00003af3ffff8e62;
    assign coff[801 ] = 64'h00003ae8ffff8e5c;
    assign coff[802 ] = 64'h00003addffff8e56;
    assign coff[803 ] = 64'h00003ad1ffff8e50;
    assign coff[804 ] = 64'h00003ac6ffff8e4b;
    assign coff[805 ] = 64'h00003abbffff8e45;
    assign coff[806 ] = 64'h00003ab0ffff8e3f;
    assign coff[807 ] = 64'h00003aa5ffff8e39;
    assign coff[808 ] = 64'h00003a9affff8e34;
    assign coff[809 ] = 64'h00003a8effff8e2e;
    assign coff[810 ] = 64'h00003a83ffff8e28;
    assign coff[811 ] = 64'h00003a78ffff8e22;
    assign coff[812 ] = 64'h00003a6dffff8e1d;
    assign coff[813 ] = 64'h00003a62ffff8e17;
    assign coff[814 ] = 64'h00003a57ffff8e11;
    assign coff[815 ] = 64'h00003a4bffff8e0b;
    assign coff[816 ] = 64'h00003a40ffff8e06;
    assign coff[817 ] = 64'h00003a35ffff8e00;
    assign coff[818 ] = 64'h00003a2affff8dfa;
    assign coff[819 ] = 64'h00003a1fffff8df5;
    assign coff[820 ] = 64'h00003a13ffff8def;
    assign coff[821 ] = 64'h00003a08ffff8de9;
    assign coff[822 ] = 64'h000039fdffff8de4;
    assign coff[823 ] = 64'h000039f2ffff8dde;
    assign coff[824 ] = 64'h000039e7ffff8dd8;
    assign coff[825 ] = 64'h000039dbffff8dd2;
    assign coff[826 ] = 64'h000039d0ffff8dcd;
    assign coff[827 ] = 64'h000039c5ffff8dc7;
    assign coff[828 ] = 64'h000039baffff8dc1;
    assign coff[829 ] = 64'h000039afffff8dbc;
    assign coff[830 ] = 64'h000039a3ffff8db6;
    assign coff[831 ] = 64'h00003998ffff8db0;
    assign coff[832 ] = 64'h0000398dffff8dab;
    assign coff[833 ] = 64'h00003982ffff8da5;
    assign coff[834 ] = 64'h00003976ffff8da0;
    assign coff[835 ] = 64'h0000396bffff8d9a;
    assign coff[836 ] = 64'h00003960ffff8d94;
    assign coff[837 ] = 64'h00003955ffff8d8f;
    assign coff[838 ] = 64'h00003949ffff8d89;
    assign coff[839 ] = 64'h0000393effff8d83;
    assign coff[840 ] = 64'h00003933ffff8d7e;
    assign coff[841 ] = 64'h00003928ffff8d78;
    assign coff[842 ] = 64'h0000391dffff8d73;
    assign coff[843 ] = 64'h00003911ffff8d6d;
    assign coff[844 ] = 64'h00003906ffff8d67;
    assign coff[845 ] = 64'h000038fbffff8d62;
    assign coff[846 ] = 64'h000038f0ffff8d5c;
    assign coff[847 ] = 64'h000038e4ffff8d57;
    assign coff[848 ] = 64'h000038d9ffff8d51;
    assign coff[849 ] = 64'h000038ceffff8d4b;
    assign coff[850 ] = 64'h000038c2ffff8d46;
    assign coff[851 ] = 64'h000038b7ffff8d40;
    assign coff[852 ] = 64'h000038acffff8d3b;
    assign coff[853 ] = 64'h000038a1ffff8d35;
    assign coff[854 ] = 64'h00003895ffff8d30;
    assign coff[855 ] = 64'h0000388affff8d2a;
    assign coff[856 ] = 64'h0000387fffff8d24;
    assign coff[857 ] = 64'h00003874ffff8d1f;
    assign coff[858 ] = 64'h00003868ffff8d19;
    assign coff[859 ] = 64'h0000385dffff8d14;
    assign coff[860 ] = 64'h00003852ffff8d0e;
    assign coff[861 ] = 64'h00003846ffff8d09;
    assign coff[862 ] = 64'h0000383bffff8d03;
    assign coff[863 ] = 64'h00003830ffff8cfe;
    assign coff[864 ] = 64'h00003825ffff8cf8;
    assign coff[865 ] = 64'h00003819ffff8cf3;
    assign coff[866 ] = 64'h0000380effff8ced;
    assign coff[867 ] = 64'h00003803ffff8ce8;
    assign coff[868 ] = 64'h000037f7ffff8ce2;
    assign coff[869 ] = 64'h000037ecffff8cdd;
    assign coff[870 ] = 64'h000037e1ffff8cd7;
    assign coff[871 ] = 64'h000037d5ffff8cd2;
    assign coff[872 ] = 64'h000037caffff8ccc;
    assign coff[873 ] = 64'h000037bfffff8cc7;
    assign coff[874 ] = 64'h000037b4ffff8cc1;
    assign coff[875 ] = 64'h000037a8ffff8cbc;
    assign coff[876 ] = 64'h0000379dffff8cb6;
    assign coff[877 ] = 64'h00003792ffff8cb1;
    assign coff[878 ] = 64'h00003786ffff8cab;
    assign coff[879 ] = 64'h0000377bffff8ca6;
    assign coff[880 ] = 64'h00003770ffff8ca1;
    assign coff[881 ] = 64'h00003764ffff8c9b;
    assign coff[882 ] = 64'h00003759ffff8c96;
    assign coff[883 ] = 64'h0000374effff8c90;
    assign coff[884 ] = 64'h00003742ffff8c8b;
    assign coff[885 ] = 64'h00003737ffff8c85;
    assign coff[886 ] = 64'h0000372cffff8c80;
    assign coff[887 ] = 64'h00003720ffff8c7b;
    assign coff[888 ] = 64'h00003715ffff8c75;
    assign coff[889 ] = 64'h0000370affff8c70;
    assign coff[890 ] = 64'h000036feffff8c6a;
    assign coff[891 ] = 64'h000036f3ffff8c65;
    assign coff[892 ] = 64'h000036e8ffff8c60;
    assign coff[893 ] = 64'h000036dcffff8c5a;
    assign coff[894 ] = 64'h000036d1ffff8c55;
    assign coff[895 ] = 64'h000036c5ffff8c4f;
    assign coff[896 ] = 64'h000036baffff8c4a;
    assign coff[897 ] = 64'h000036afffff8c45;
    assign coff[898 ] = 64'h000036a3ffff8c3f;
    assign coff[899 ] = 64'h00003698ffff8c3a;
    assign coff[900 ] = 64'h0000368dffff8c35;
    assign coff[901 ] = 64'h00003681ffff8c2f;
    assign coff[902 ] = 64'h00003676ffff8c2a;
    assign coff[903 ] = 64'h0000366bffff8c25;
    assign coff[904 ] = 64'h0000365fffff8c1f;
    assign coff[905 ] = 64'h00003654ffff8c1a;
    assign coff[906 ] = 64'h00003648ffff8c15;
    assign coff[907 ] = 64'h0000363dffff8c0f;
    assign coff[908 ] = 64'h00003632ffff8c0a;
    assign coff[909 ] = 64'h00003626ffff8c05;
    assign coff[910 ] = 64'h0000361bffff8bff;
    assign coff[911 ] = 64'h0000360fffff8bfa;
    assign coff[912 ] = 64'h00003604ffff8bf5;
    assign coff[913 ] = 64'h000035f9ffff8bef;
    assign coff[914 ] = 64'h000035edffff8bea;
    assign coff[915 ] = 64'h000035e2ffff8be5;
    assign coff[916 ] = 64'h000035d7ffff8bdf;
    assign coff[917 ] = 64'h000035cbffff8bda;
    assign coff[918 ] = 64'h000035c0ffff8bd5;
    assign coff[919 ] = 64'h000035b4ffff8bd0;
    assign coff[920 ] = 64'h000035a9ffff8bca;
    assign coff[921 ] = 64'h0000359dffff8bc5;
    assign coff[922 ] = 64'h00003592ffff8bc0;
    assign coff[923 ] = 64'h00003587ffff8bbb;
    assign coff[924 ] = 64'h0000357bffff8bb5;
    assign coff[925 ] = 64'h00003570ffff8bb0;
    assign coff[926 ] = 64'h00003564ffff8bab;
    assign coff[927 ] = 64'h00003559ffff8ba6;
    assign coff[928 ] = 64'h0000354effff8ba0;
    assign coff[929 ] = 64'h00003542ffff8b9b;
    assign coff[930 ] = 64'h00003537ffff8b96;
    assign coff[931 ] = 64'h0000352bffff8b91;
    assign coff[932 ] = 64'h00003520ffff8b8b;
    assign coff[933 ] = 64'h00003514ffff8b86;
    assign coff[934 ] = 64'h00003509ffff8b81;
    assign coff[935 ] = 64'h000034feffff8b7c;
    assign coff[936 ] = 64'h000034f2ffff8b77;
    assign coff[937 ] = 64'h000034e7ffff8b71;
    assign coff[938 ] = 64'h000034dbffff8b6c;
    assign coff[939 ] = 64'h000034d0ffff8b67;
    assign coff[940 ] = 64'h000034c4ffff8b62;
    assign coff[941 ] = 64'h000034b9ffff8b5d;
    assign coff[942 ] = 64'h000034adffff8b58;
    assign coff[943 ] = 64'h000034a2ffff8b52;
    assign coff[944 ] = 64'h00003497ffff8b4d;
    assign coff[945 ] = 64'h0000348bffff8b48;
    assign coff[946 ] = 64'h00003480ffff8b43;
    assign coff[947 ] = 64'h00003474ffff8b3e;
    assign coff[948 ] = 64'h00003469ffff8b39;
    assign coff[949 ] = 64'h0000345dffff8b33;
    assign coff[950 ] = 64'h00003452ffff8b2e;
    assign coff[951 ] = 64'h00003446ffff8b29;
    assign coff[952 ] = 64'h0000343bffff8b24;
    assign coff[953 ] = 64'h0000342fffff8b1f;
    assign coff[954 ] = 64'h00003424ffff8b1a;
    assign coff[955 ] = 64'h00003418ffff8b15;
    assign coff[956 ] = 64'h0000340dffff8b10;
    assign coff[957 ] = 64'h00003401ffff8b0a;
    assign coff[958 ] = 64'h000033f6ffff8b05;
    assign coff[959 ] = 64'h000033eaffff8b00;
    assign coff[960 ] = 64'h000033dfffff8afb;
    assign coff[961 ] = 64'h000033d3ffff8af6;
    assign coff[962 ] = 64'h000033c8ffff8af1;
    assign coff[963 ] = 64'h000033bcffff8aec;
    assign coff[964 ] = 64'h000033b1ffff8ae7;
    assign coff[965 ] = 64'h000033a5ffff8ae2;
    assign coff[966 ] = 64'h0000339affff8add;
    assign coff[967 ] = 64'h0000338effff8ad8;
    assign coff[968 ] = 64'h00003383ffff8ad3;
    assign coff[969 ] = 64'h00003377ffff8ace;
    assign coff[970 ] = 64'h0000336cffff8ac8;
    assign coff[971 ] = 64'h00003360ffff8ac3;
    assign coff[972 ] = 64'h00003355ffff8abe;
    assign coff[973 ] = 64'h00003349ffff8ab9;
    assign coff[974 ] = 64'h0000333effff8ab4;
    assign coff[975 ] = 64'h00003332ffff8aaf;
    assign coff[976 ] = 64'h00003327ffff8aaa;
    assign coff[977 ] = 64'h0000331bffff8aa5;
    assign coff[978 ] = 64'h00003310ffff8aa0;
    assign coff[979 ] = 64'h00003304ffff8a9b;
    assign coff[980 ] = 64'h000032f9ffff8a96;
    assign coff[981 ] = 64'h000032edffff8a91;
    assign coff[982 ] = 64'h000032e2ffff8a8c;
    assign coff[983 ] = 64'h000032d6ffff8a87;
    assign coff[984 ] = 64'h000032cbffff8a82;
    assign coff[985 ] = 64'h000032bfffff8a7d;
    assign coff[986 ] = 64'h000032b4ffff8a78;
    assign coff[987 ] = 64'h000032a8ffff8a73;
    assign coff[988 ] = 64'h0000329dffff8a6e;
    assign coff[989 ] = 64'h00003291ffff8a69;
    assign coff[990 ] = 64'h00003285ffff8a64;
    assign coff[991 ] = 64'h0000327affff8a5f;
    assign coff[992 ] = 64'h0000326effff8a5a;
    assign coff[993 ] = 64'h00003263ffff8a56;
    assign coff[994 ] = 64'h00003257ffff8a51;
    assign coff[995 ] = 64'h0000324cffff8a4c;
    assign coff[996 ] = 64'h00003240ffff8a47;
    assign coff[997 ] = 64'h00003235ffff8a42;
    assign coff[998 ] = 64'h00003229ffff8a3d;
    assign coff[999 ] = 64'h0000321dffff8a38;
    assign coff[1000] = 64'h00003212ffff8a33;
    assign coff[1001] = 64'h00003206ffff8a2e;
    assign coff[1002] = 64'h000031fbffff8a29;
    assign coff[1003] = 64'h000031efffff8a24;
    assign coff[1004] = 64'h000031e4ffff8a1f;
    assign coff[1005] = 64'h000031d8ffff8a1a;
    assign coff[1006] = 64'h000031ccffff8a16;
    assign coff[1007] = 64'h000031c1ffff8a11;
    assign coff[1008] = 64'h000031b5ffff8a0c;
    assign coff[1009] = 64'h000031aaffff8a07;
    assign coff[1010] = 64'h0000319effff8a02;
    assign coff[1011] = 64'h00003193ffff89fd;
    assign coff[1012] = 64'h00003187ffff89f8;
    assign coff[1013] = 64'h0000317bffff89f3;
    assign coff[1014] = 64'h00003170ffff89ef;
    assign coff[1015] = 64'h00003164ffff89ea;
    assign coff[1016] = 64'h00003159ffff89e5;
    assign coff[1017] = 64'h0000314dffff89e0;
    assign coff[1018] = 64'h00003141ffff89db;
    assign coff[1019] = 64'h00003136ffff89d6;
    assign coff[1020] = 64'h0000312affff89d2;
    assign coff[1021] = 64'h0000311fffff89cd;
    assign coff[1022] = 64'h00003113ffff89c8;
    assign coff[1023] = 64'h00003107ffff89c3;
    assign coff[1024] = 64'h000030fcffff89be;
    assign coff[1025] = 64'h000030f0ffff89ba;
    assign coff[1026] = 64'h000030e5ffff89b5;
    assign coff[1027] = 64'h000030d9ffff89b0;
    assign coff[1028] = 64'h000030cdffff89ab;
    assign coff[1029] = 64'h000030c2ffff89a6;
    assign coff[1030] = 64'h000030b6ffff89a2;
    assign coff[1031] = 64'h000030aaffff899d;
    assign coff[1032] = 64'h0000309fffff8998;
    assign coff[1033] = 64'h00003093ffff8993;
    assign coff[1034] = 64'h00003088ffff898e;
    assign coff[1035] = 64'h0000307cffff898a;
    assign coff[1036] = 64'h00003070ffff8985;
    assign coff[1037] = 64'h00003065ffff8980;
    assign coff[1038] = 64'h00003059ffff897b;
    assign coff[1039] = 64'h0000304dffff8977;
    assign coff[1040] = 64'h00003042ffff8972;
    assign coff[1041] = 64'h00003036ffff896d;
    assign coff[1042] = 64'h0000302affff8968;
    assign coff[1043] = 64'h0000301fffff8964;
    assign coff[1044] = 64'h00003013ffff895f;
    assign coff[1045] = 64'h00003008ffff895a;
    assign coff[1046] = 64'h00002ffcffff8956;
    assign coff[1047] = 64'h00002ff0ffff8951;
    assign coff[1048] = 64'h00002fe5ffff894c;
    assign coff[1049] = 64'h00002fd9ffff8947;
    assign coff[1050] = 64'h00002fcdffff8943;
    assign coff[1051] = 64'h00002fc2ffff893e;
    assign coff[1052] = 64'h00002fb6ffff8939;
    assign coff[1053] = 64'h00002faaffff8935;
    assign coff[1054] = 64'h00002f9fffff8930;
    assign coff[1055] = 64'h00002f93ffff892b;
    assign coff[1056] = 64'h00002f87ffff8927;
    assign coff[1057] = 64'h00002f7cffff8922;
    assign coff[1058] = 64'h00002f70ffff891d;
    assign coff[1059] = 64'h00002f64ffff8919;
    assign coff[1060] = 64'h00002f59ffff8914;
    assign coff[1061] = 64'h00002f4dffff890f;
    assign coff[1062] = 64'h00002f41ffff890b;
    assign coff[1063] = 64'h00002f36ffff8906;
    assign coff[1064] = 64'h00002f2affff8902;
    assign coff[1065] = 64'h00002f1effff88fd;
    assign coff[1066] = 64'h00002f13ffff88f8;
    assign coff[1067] = 64'h00002f07ffff88f4;
    assign coff[1068] = 64'h00002efbffff88ef;
    assign coff[1069] = 64'h00002eefffff88ea;
    assign coff[1070] = 64'h00002ee4ffff88e6;
    assign coff[1071] = 64'h00002ed8ffff88e1;
    assign coff[1072] = 64'h00002eccffff88dd;
    assign coff[1073] = 64'h00002ec1ffff88d8;
    assign coff[1074] = 64'h00002eb5ffff88d3;
    assign coff[1075] = 64'h00002ea9ffff88cf;
    assign coff[1076] = 64'h00002e9effff88ca;
    assign coff[1077] = 64'h00002e92ffff88c6;
    assign coff[1078] = 64'h00002e86ffff88c1;
    assign coff[1079] = 64'h00002e7affff88bd;
    assign coff[1080] = 64'h00002e6fffff88b8;
    assign coff[1081] = 64'h00002e63ffff88b3;
    assign coff[1082] = 64'h00002e57ffff88af;
    assign coff[1083] = 64'h00002e4cffff88aa;
    assign coff[1084] = 64'h00002e40ffff88a6;
    assign coff[1085] = 64'h00002e34ffff88a1;
    assign coff[1086] = 64'h00002e28ffff889d;
    assign coff[1087] = 64'h00002e1dffff8898;
    assign coff[1088] = 64'h00002e11ffff8894;
    assign coff[1089] = 64'h00002e05ffff888f;
    assign coff[1090] = 64'h00002dfaffff888b;
    assign coff[1091] = 64'h00002deeffff8886;
    assign coff[1092] = 64'h00002de2ffff8882;
    assign coff[1093] = 64'h00002dd6ffff887d;
    assign coff[1094] = 64'h00002dcbffff8879;
    assign coff[1095] = 64'h00002dbfffff8874;
    assign coff[1096] = 64'h00002db3ffff8870;
    assign coff[1097] = 64'h00002da7ffff886b;
    assign coff[1098] = 64'h00002d9cffff8867;
    assign coff[1099] = 64'h00002d90ffff8862;
    assign coff[1100] = 64'h00002d84ffff885e;
    assign coff[1101] = 64'h00002d78ffff8859;
    assign coff[1102] = 64'h00002d6dffff8855;
    assign coff[1103] = 64'h00002d61ffff8850;
    assign coff[1104] = 64'h00002d55ffff884c;
    assign coff[1105] = 64'h00002d49ffff8847;
    assign coff[1106] = 64'h00002d3effff8843;
    assign coff[1107] = 64'h00002d32ffff883f;
    assign coff[1108] = 64'h00002d26ffff883a;
    assign coff[1109] = 64'h00002d1affff8836;
    assign coff[1110] = 64'h00002d0fffff8831;
    assign coff[1111] = 64'h00002d03ffff882d;
    assign coff[1112] = 64'h00002cf7ffff8828;
    assign coff[1113] = 64'h00002cebffff8824;
    assign coff[1114] = 64'h00002ce0ffff8820;
    assign coff[1115] = 64'h00002cd4ffff881b;
    assign coff[1116] = 64'h00002cc8ffff8817;
    assign coff[1117] = 64'h00002cbcffff8812;
    assign coff[1118] = 64'h00002cb1ffff880e;
    assign coff[1119] = 64'h00002ca5ffff880a;
    assign coff[1120] = 64'h00002c99ffff8805;
    assign coff[1121] = 64'h00002c8dffff8801;
    assign coff[1122] = 64'h00002c81ffff87fd;
    assign coff[1123] = 64'h00002c76ffff87f8;
    assign coff[1124] = 64'h00002c6affff87f4;
    assign coff[1125] = 64'h00002c5effff87ef;
    assign coff[1126] = 64'h00002c52ffff87eb;
    assign coff[1127] = 64'h00002c46ffff87e7;
    assign coff[1128] = 64'h00002c3bffff87e2;
    assign coff[1129] = 64'h00002c2fffff87de;
    assign coff[1130] = 64'h00002c23ffff87da;
    assign coff[1131] = 64'h00002c17ffff87d5;
    assign coff[1132] = 64'h00002c0cffff87d1;
    assign coff[1133] = 64'h00002c00ffff87cd;
    assign coff[1134] = 64'h00002bf4ffff87c8;
    assign coff[1135] = 64'h00002be8ffff87c4;
    assign coff[1136] = 64'h00002bdcffff87c0;
    assign coff[1137] = 64'h00002bd0ffff87bb;
    assign coff[1138] = 64'h00002bc5ffff87b7;
    assign coff[1139] = 64'h00002bb9ffff87b3;
    assign coff[1140] = 64'h00002badffff87af;
    assign coff[1141] = 64'h00002ba1ffff87aa;
    assign coff[1142] = 64'h00002b95ffff87a6;
    assign coff[1143] = 64'h00002b8affff87a2;
    assign coff[1144] = 64'h00002b7effff879d;
    assign coff[1145] = 64'h00002b72ffff8799;
    assign coff[1146] = 64'h00002b66ffff8795;
    assign coff[1147] = 64'h00002b5affff8791;
    assign coff[1148] = 64'h00002b4fffff878c;
    assign coff[1149] = 64'h00002b43ffff8788;
    assign coff[1150] = 64'h00002b37ffff8784;
    assign coff[1151] = 64'h00002b2bffff8780;
    assign coff[1152] = 64'h00002b1fffff877b;
    assign coff[1153] = 64'h00002b13ffff8777;
    assign coff[1154] = 64'h00002b08ffff8773;
    assign coff[1155] = 64'h00002afcffff876f;
    assign coff[1156] = 64'h00002af0ffff876b;
    assign coff[1157] = 64'h00002ae4ffff8766;
    assign coff[1158] = 64'h00002ad8ffff8762;
    assign coff[1159] = 64'h00002accffff875e;
    assign coff[1160] = 64'h00002ac1ffff875a;
    assign coff[1161] = 64'h00002ab5ffff8756;
    assign coff[1162] = 64'h00002aa9ffff8751;
    assign coff[1163] = 64'h00002a9dffff874d;
    assign coff[1164] = 64'h00002a91ffff8749;
    assign coff[1165] = 64'h00002a85ffff8745;
    assign coff[1166] = 64'h00002a79ffff8741;
    assign coff[1167] = 64'h00002a6effff873c;
    assign coff[1168] = 64'h00002a62ffff8738;
    assign coff[1169] = 64'h00002a56ffff8734;
    assign coff[1170] = 64'h00002a4affff8730;
    assign coff[1171] = 64'h00002a3effff872c;
    assign coff[1172] = 64'h00002a32ffff8728;
    assign coff[1173] = 64'h00002a26ffff8724;
    assign coff[1174] = 64'h00002a1bffff871f;
    assign coff[1175] = 64'h00002a0fffff871b;
    assign coff[1176] = 64'h00002a03ffff8717;
    assign coff[1177] = 64'h000029f7ffff8713;
    assign coff[1178] = 64'h000029ebffff870f;
    assign coff[1179] = 64'h000029dfffff870b;
    assign coff[1180] = 64'h000029d3ffff8707;
    assign coff[1181] = 64'h000029c7ffff8703;
    assign coff[1182] = 64'h000029bcffff86ff;
    assign coff[1183] = 64'h000029b0ffff86fa;
    assign coff[1184] = 64'h000029a4ffff86f6;
    assign coff[1185] = 64'h00002998ffff86f2;
    assign coff[1186] = 64'h0000298cffff86ee;
    assign coff[1187] = 64'h00002980ffff86ea;
    assign coff[1188] = 64'h00002974ffff86e6;
    assign coff[1189] = 64'h00002968ffff86e2;
    assign coff[1190] = 64'h0000295cffff86de;
    assign coff[1191] = 64'h00002951ffff86da;
    assign coff[1192] = 64'h00002945ffff86d6;
    assign coff[1193] = 64'h00002939ffff86d2;
    assign coff[1194] = 64'h0000292dffff86ce;
    assign coff[1195] = 64'h00002921ffff86ca;
    assign coff[1196] = 64'h00002915ffff86c6;
    assign coff[1197] = 64'h00002909ffff86c2;
    assign coff[1198] = 64'h000028fdffff86be;
    assign coff[1199] = 64'h000028f1ffff86ba;
    assign coff[1200] = 64'h000028e5ffff86b6;
    assign coff[1201] = 64'h000028daffff86b2;
    assign coff[1202] = 64'h000028ceffff86ad;
    assign coff[1203] = 64'h000028c2ffff86a9;
    assign coff[1204] = 64'h000028b6ffff86a5;
    assign coff[1205] = 64'h000028aaffff86a1;
    assign coff[1206] = 64'h0000289effff869e;
    assign coff[1207] = 64'h00002892ffff869a;
    assign coff[1208] = 64'h00002886ffff8696;
    assign coff[1209] = 64'h0000287affff8692;
    assign coff[1210] = 64'h0000286effff868e;
    assign coff[1211] = 64'h00002862ffff868a;
    assign coff[1212] = 64'h00002856ffff8686;
    assign coff[1213] = 64'h0000284bffff8682;
    assign coff[1214] = 64'h0000283fffff867e;
    assign coff[1215] = 64'h00002833ffff867a;
    assign coff[1216] = 64'h00002827ffff8676;
    assign coff[1217] = 64'h0000281bffff8672;
    assign coff[1218] = 64'h0000280fffff866e;
    assign coff[1219] = 64'h00002803ffff866a;
    assign coff[1220] = 64'h000027f7ffff8666;
    assign coff[1221] = 64'h000027ebffff8662;
    assign coff[1222] = 64'h000027dfffff865e;
    assign coff[1223] = 64'h000027d3ffff865a;
    assign coff[1224] = 64'h000027c7ffff8656;
    assign coff[1225] = 64'h000027bbffff8653;
    assign coff[1226] = 64'h000027afffff864f;
    assign coff[1227] = 64'h000027a3ffff864b;
    assign coff[1228] = 64'h00002797ffff8647;
    assign coff[1229] = 64'h0000278bffff8643;
    assign coff[1230] = 64'h00002780ffff863f;
    assign coff[1231] = 64'h00002774ffff863b;
    assign coff[1232] = 64'h00002768ffff8637;
    assign coff[1233] = 64'h0000275cffff8634;
    assign coff[1234] = 64'h00002750ffff8630;
    assign coff[1235] = 64'h00002744ffff862c;
    assign coff[1236] = 64'h00002738ffff8628;
    assign coff[1237] = 64'h0000272cffff8624;
    assign coff[1238] = 64'h00002720ffff8620;
    assign coff[1239] = 64'h00002714ffff861c;
    assign coff[1240] = 64'h00002708ffff8619;
    assign coff[1241] = 64'h000026fcffff8615;
    assign coff[1242] = 64'h000026f0ffff8611;
    assign coff[1243] = 64'h000026e4ffff860d;
    assign coff[1244] = 64'h000026d8ffff8609;
    assign coff[1245] = 64'h000026ccffff8605;
    assign coff[1246] = 64'h000026c0ffff8602;
    assign coff[1247] = 64'h000026b4ffff85fe;
    assign coff[1248] = 64'h000026a8ffff85fa;
    assign coff[1249] = 64'h0000269cffff85f6;
    assign coff[1250] = 64'h00002690ffff85f2;
    assign coff[1251] = 64'h00002684ffff85ef;
    assign coff[1252] = 64'h00002678ffff85eb;
    assign coff[1253] = 64'h0000266cffff85e7;
    assign coff[1254] = 64'h00002660ffff85e3;
    assign coff[1255] = 64'h00002654ffff85e0;
    assign coff[1256] = 64'h00002648ffff85dc;
    assign coff[1257] = 64'h0000263cffff85d8;
    assign coff[1258] = 64'h00002630ffff85d4;
    assign coff[1259] = 64'h00002624ffff85d1;
    assign coff[1260] = 64'h00002618ffff85cd;
    assign coff[1261] = 64'h0000260cffff85c9;
    assign coff[1262] = 64'h00002600ffff85c5;
    assign coff[1263] = 64'h000025f4ffff85c2;
    assign coff[1264] = 64'h000025e8ffff85be;
    assign coff[1265] = 64'h000025dcffff85ba;
    assign coff[1266] = 64'h000025d0ffff85b7;
    assign coff[1267] = 64'h000025c4ffff85b3;
    assign coff[1268] = 64'h000025b8ffff85af;
    assign coff[1269] = 64'h000025acffff85ab;
    assign coff[1270] = 64'h000025a0ffff85a8;
    assign coff[1271] = 64'h00002594ffff85a4;
    assign coff[1272] = 64'h00002588ffff85a0;
    assign coff[1273] = 64'h0000257cffff859d;
    assign coff[1274] = 64'h00002570ffff8599;
    assign coff[1275] = 64'h00002564ffff8595;
    assign coff[1276] = 64'h00002558ffff8592;
    assign coff[1277] = 64'h0000254cffff858e;
    assign coff[1278] = 64'h00002540ffff858a;
    assign coff[1279] = 64'h00002534ffff8587;
    assign coff[1280] = 64'h00002528ffff8583;
    assign coff[1281] = 64'h0000251cffff857f;
    assign coff[1282] = 64'h00002510ffff857c;
    assign coff[1283] = 64'h00002504ffff8578;
    assign coff[1284] = 64'h000024f8ffff8574;
    assign coff[1285] = 64'h000024ecffff8571;
    assign coff[1286] = 64'h000024e0ffff856d;
    assign coff[1287] = 64'h000024d4ffff856a;
    assign coff[1288] = 64'h000024c8ffff8566;
    assign coff[1289] = 64'h000024bcffff8562;
    assign coff[1290] = 64'h000024b0ffff855f;
    assign coff[1291] = 64'h000024a4ffff855b;
    assign coff[1292] = 64'h00002498ffff8558;
    assign coff[1293] = 64'h0000248cffff8554;
    assign coff[1294] = 64'h00002480ffff8550;
    assign coff[1295] = 64'h00002474ffff854d;
    assign coff[1296] = 64'h00002467ffff8549;
    assign coff[1297] = 64'h0000245bffff8546;
    assign coff[1298] = 64'h0000244fffff8542;
    assign coff[1299] = 64'h00002443ffff853f;
    assign coff[1300] = 64'h00002437ffff853b;
    assign coff[1301] = 64'h0000242bffff8537;
    assign coff[1302] = 64'h0000241fffff8534;
    assign coff[1303] = 64'h00002413ffff8530;
    assign coff[1304] = 64'h00002407ffff852d;
    assign coff[1305] = 64'h000023fbffff8529;
    assign coff[1306] = 64'h000023efffff8526;
    assign coff[1307] = 64'h000023e3ffff8522;
    assign coff[1308] = 64'h000023d7ffff851f;
    assign coff[1309] = 64'h000023cbffff851b;
    assign coff[1310] = 64'h000023bfffff8518;
    assign coff[1311] = 64'h000023b3ffff8514;
    assign coff[1312] = 64'h000023a7ffff8511;
    assign coff[1313] = 64'h0000239affff850d;
    assign coff[1314] = 64'h0000238effff850a;
    assign coff[1315] = 64'h00002382ffff8506;
    assign coff[1316] = 64'h00002376ffff8503;
    assign coff[1317] = 64'h0000236affff84ff;
    assign coff[1318] = 64'h0000235effff84fc;
    assign coff[1319] = 64'h00002352ffff84f8;
    assign coff[1320] = 64'h00002346ffff84f5;
    assign coff[1321] = 64'h0000233affff84f1;
    assign coff[1322] = 64'h0000232effff84ee;
    assign coff[1323] = 64'h00002322ffff84ea;
    assign coff[1324] = 64'h00002316ffff84e7;
    assign coff[1325] = 64'h0000230affff84e4;
    assign coff[1326] = 64'h000022fdffff84e0;
    assign coff[1327] = 64'h000022f1ffff84dd;
    assign coff[1328] = 64'h000022e5ffff84d9;
    assign coff[1329] = 64'h000022d9ffff84d6;
    assign coff[1330] = 64'h000022cdffff84d2;
    assign coff[1331] = 64'h000022c1ffff84cf;
    assign coff[1332] = 64'h000022b5ffff84cc;
    assign coff[1333] = 64'h000022a9ffff84c8;
    assign coff[1334] = 64'h0000229dffff84c5;
    assign coff[1335] = 64'h00002291ffff84c1;
    assign coff[1336] = 64'h00002284ffff84be;
    assign coff[1337] = 64'h00002278ffff84bb;
    assign coff[1338] = 64'h0000226cffff84b7;
    assign coff[1339] = 64'h00002260ffff84b4;
    assign coff[1340] = 64'h00002254ffff84b0;
    assign coff[1341] = 64'h00002248ffff84ad;
    assign coff[1342] = 64'h0000223cffff84aa;
    assign coff[1343] = 64'h00002230ffff84a6;
    assign coff[1344] = 64'h00002224ffff84a3;
    assign coff[1345] = 64'h00002218ffff84a0;
    assign coff[1346] = 64'h0000220bffff849c;
    assign coff[1347] = 64'h000021ffffff8499;
    assign coff[1348] = 64'h000021f3ffff8496;
    assign coff[1349] = 64'h000021e7ffff8492;
    assign coff[1350] = 64'h000021dbffff848f;
    assign coff[1351] = 64'h000021cfffff848c;
    assign coff[1352] = 64'h000021c3ffff8488;
    assign coff[1353] = 64'h000021b7ffff8485;
    assign coff[1354] = 64'h000021aaffff8482;
    assign coff[1355] = 64'h0000219effff847e;
    assign coff[1356] = 64'h00002192ffff847b;
    assign coff[1357] = 64'h00002186ffff8478;
    assign coff[1358] = 64'h0000217affff8475;
    assign coff[1359] = 64'h0000216effff8471;
    assign coff[1360] = 64'h00002162ffff846e;
    assign coff[1361] = 64'h00002156ffff846b;
    assign coff[1362] = 64'h00002149ffff8467;
    assign coff[1363] = 64'h0000213dffff8464;
    assign coff[1364] = 64'h00002131ffff8461;
    assign coff[1365] = 64'h00002125ffff845e;
    assign coff[1366] = 64'h00002119ffff845a;
    assign coff[1367] = 64'h0000210dffff8457;
    assign coff[1368] = 64'h00002101ffff8454;
    assign coff[1369] = 64'h000020f4ffff8451;
    assign coff[1370] = 64'h000020e8ffff844d;
    assign coff[1371] = 64'h000020dcffff844a;
    assign coff[1372] = 64'h000020d0ffff8447;
    assign coff[1373] = 64'h000020c4ffff8444;
    assign coff[1374] = 64'h000020b8ffff8441;
    assign coff[1375] = 64'h000020acffff843d;
    assign coff[1376] = 64'h0000209fffff843a;
    assign coff[1377] = 64'h00002093ffff8437;
    assign coff[1378] = 64'h00002087ffff8434;
    assign coff[1379] = 64'h0000207bffff8431;
    assign coff[1380] = 64'h0000206fffff842d;
    assign coff[1381] = 64'h00002063ffff842a;
    assign coff[1382] = 64'h00002057ffff8427;
    assign coff[1383] = 64'h0000204affff8424;
    assign coff[1384] = 64'h0000203effff8421;
    assign coff[1385] = 64'h00002032ffff841d;
    assign coff[1386] = 64'h00002026ffff841a;
    assign coff[1387] = 64'h0000201affff8417;
    assign coff[1388] = 64'h0000200effff8414;
    assign coff[1389] = 64'h00002001ffff8411;
    assign coff[1390] = 64'h00001ff5ffff840e;
    assign coff[1391] = 64'h00001fe9ffff840b;
    assign coff[1392] = 64'h00001fddffff8407;
    assign coff[1393] = 64'h00001fd1ffff8404;
    assign coff[1394] = 64'h00001fc5ffff8401;
    assign coff[1395] = 64'h00001fb8ffff83fe;
    assign coff[1396] = 64'h00001facffff83fb;
    assign coff[1397] = 64'h00001fa0ffff83f8;
    assign coff[1398] = 64'h00001f94ffff83f5;
    assign coff[1399] = 64'h00001f88ffff83f2;
    assign coff[1400] = 64'h00001f7bffff83ef;
    assign coff[1401] = 64'h00001f6fffff83ec;
    assign coff[1402] = 64'h00001f63ffff83e8;
    assign coff[1403] = 64'h00001f57ffff83e5;
    assign coff[1404] = 64'h00001f4bffff83e2;
    assign coff[1405] = 64'h00001f3fffff83df;
    assign coff[1406] = 64'h00001f32ffff83dc;
    assign coff[1407] = 64'h00001f26ffff83d9;
    assign coff[1408] = 64'h00001f1affff83d6;
    assign coff[1409] = 64'h00001f0effff83d3;
    assign coff[1410] = 64'h00001f02ffff83d0;
    assign coff[1411] = 64'h00001ef5ffff83cd;
    assign coff[1412] = 64'h00001ee9ffff83ca;
    assign coff[1413] = 64'h00001eddffff83c7;
    assign coff[1414] = 64'h00001ed1ffff83c4;
    assign coff[1415] = 64'h00001ec5ffff83c1;
    assign coff[1416] = 64'h00001eb8ffff83be;
    assign coff[1417] = 64'h00001eacffff83bb;
    assign coff[1418] = 64'h00001ea0ffff83b8;
    assign coff[1419] = 64'h00001e94ffff83b5;
    assign coff[1420] = 64'h00001e88ffff83b2;
    assign coff[1421] = 64'h00001e7bffff83af;
    assign coff[1422] = 64'h00001e6fffff83ac;
    assign coff[1423] = 64'h00001e63ffff83a9;
    assign coff[1424] = 64'h00001e57ffff83a6;
    assign coff[1425] = 64'h00001e4bffff83a3;
    assign coff[1426] = 64'h00001e3effff83a0;
    assign coff[1427] = 64'h00001e32ffff839d;
    assign coff[1428] = 64'h00001e26ffff839a;
    assign coff[1429] = 64'h00001e1affff8397;
    assign coff[1430] = 64'h00001e0effff8394;
    assign coff[1431] = 64'h00001e01ffff8391;
    assign coff[1432] = 64'h00001df5ffff838e;
    assign coff[1433] = 64'h00001de9ffff838b;
    assign coff[1434] = 64'h00001dddffff8388;
    assign coff[1435] = 64'h00001dd0ffff8385;
    assign coff[1436] = 64'h00001dc4ffff8382;
    assign coff[1437] = 64'h00001db8ffff837f;
    assign coff[1438] = 64'h00001dacffff837d;
    assign coff[1439] = 64'h00001da0ffff837a;
    assign coff[1440] = 64'h00001d93ffff8377;
    assign coff[1441] = 64'h00001d87ffff8374;
    assign coff[1442] = 64'h00001d7bffff8371;
    assign coff[1443] = 64'h00001d6fffff836e;
    assign coff[1444] = 64'h00001d62ffff836b;
    assign coff[1445] = 64'h00001d56ffff8368;
    assign coff[1446] = 64'h00001d4affff8365;
    assign coff[1447] = 64'h00001d3effff8362;
    assign coff[1448] = 64'h00001d31ffff8360;
    assign coff[1449] = 64'h00001d25ffff835d;
    assign coff[1450] = 64'h00001d19ffff835a;
    assign coff[1451] = 64'h00001d0dffff8357;
    assign coff[1452] = 64'h00001d01ffff8354;
    assign coff[1453] = 64'h00001cf4ffff8351;
    assign coff[1454] = 64'h00001ce8ffff834f;
    assign coff[1455] = 64'h00001cdcffff834c;
    assign coff[1456] = 64'h00001cd0ffff8349;
    assign coff[1457] = 64'h00001cc3ffff8346;
    assign coff[1458] = 64'h00001cb7ffff8343;
    assign coff[1459] = 64'h00001cabffff8340;
    assign coff[1460] = 64'h00001c9fffff833e;
    assign coff[1461] = 64'h00001c92ffff833b;
    assign coff[1462] = 64'h00001c86ffff8338;
    assign coff[1463] = 64'h00001c7affff8335;
    assign coff[1464] = 64'h00001c6effff8332;
    assign coff[1465] = 64'h00001c61ffff8330;
    assign coff[1466] = 64'h00001c55ffff832d;
    assign coff[1467] = 64'h00001c49ffff832a;
    assign coff[1468] = 64'h00001c3dffff8327;
    assign coff[1469] = 64'h00001c30ffff8324;
    assign coff[1470] = 64'h00001c24ffff8322;
    assign coff[1471] = 64'h00001c18ffff831f;
    assign coff[1472] = 64'h00001c0cffff831c;
    assign coff[1473] = 64'h00001bffffff8319;
    assign coff[1474] = 64'h00001bf3ffff8317;
    assign coff[1475] = 64'h00001be7ffff8314;
    assign coff[1476] = 64'h00001bdaffff8311;
    assign coff[1477] = 64'h00001bceffff830e;
    assign coff[1478] = 64'h00001bc2ffff830c;
    assign coff[1479] = 64'h00001bb6ffff8309;
    assign coff[1480] = 64'h00001ba9ffff8306;
    assign coff[1481] = 64'h00001b9dffff8304;
    assign coff[1482] = 64'h00001b91ffff8301;
    assign coff[1483] = 64'h00001b85ffff82fe;
    assign coff[1484] = 64'h00001b78ffff82fb;
    assign coff[1485] = 64'h00001b6cffff82f9;
    assign coff[1486] = 64'h00001b60ffff82f6;
    assign coff[1487] = 64'h00001b53ffff82f3;
    assign coff[1488] = 64'h00001b47ffff82f1;
    assign coff[1489] = 64'h00001b3bffff82ee;
    assign coff[1490] = 64'h00001b2fffff82eb;
    assign coff[1491] = 64'h00001b22ffff82e9;
    assign coff[1492] = 64'h00001b16ffff82e6;
    assign coff[1493] = 64'h00001b0affff82e3;
    assign coff[1494] = 64'h00001afeffff82e1;
    assign coff[1495] = 64'h00001af1ffff82de;
    assign coff[1496] = 64'h00001ae5ffff82db;
    assign coff[1497] = 64'h00001ad9ffff82d9;
    assign coff[1498] = 64'h00001accffff82d6;
    assign coff[1499] = 64'h00001ac0ffff82d4;
    assign coff[1500] = 64'h00001ab4ffff82d1;
    assign coff[1501] = 64'h00001aa8ffff82ce;
    assign coff[1502] = 64'h00001a9bffff82cc;
    assign coff[1503] = 64'h00001a8fffff82c9;
    assign coff[1504] = 64'h00001a83ffff82c6;
    assign coff[1505] = 64'h00001a76ffff82c4;
    assign coff[1506] = 64'h00001a6affff82c1;
    assign coff[1507] = 64'h00001a5effff82bf;
    assign coff[1508] = 64'h00001a51ffff82bc;
    assign coff[1509] = 64'h00001a45ffff82ba;
    assign coff[1510] = 64'h00001a39ffff82b7;
    assign coff[1511] = 64'h00001a2dffff82b4;
    assign coff[1512] = 64'h00001a20ffff82b2;
    assign coff[1513] = 64'h00001a14ffff82af;
    assign coff[1514] = 64'h00001a08ffff82ad;
    assign coff[1515] = 64'h000019fbffff82aa;
    assign coff[1516] = 64'h000019efffff82a8;
    assign coff[1517] = 64'h000019e3ffff82a5;
    assign coff[1518] = 64'h000019d6ffff82a3;
    assign coff[1519] = 64'h000019caffff82a0;
    assign coff[1520] = 64'h000019beffff829d;
    assign coff[1521] = 64'h000019b1ffff829b;
    assign coff[1522] = 64'h000019a5ffff8298;
    assign coff[1523] = 64'h00001999ffff8296;
    assign coff[1524] = 64'h0000198dffff8293;
    assign coff[1525] = 64'h00001980ffff8291;
    assign coff[1526] = 64'h00001974ffff828e;
    assign coff[1527] = 64'h00001968ffff828c;
    assign coff[1528] = 64'h0000195bffff8289;
    assign coff[1529] = 64'h0000194fffff8287;
    assign coff[1530] = 64'h00001943ffff8284;
    assign coff[1531] = 64'h00001936ffff8282;
    assign coff[1532] = 64'h0000192affff827f;
    assign coff[1533] = 64'h0000191effff827d;
    assign coff[1534] = 64'h00001911ffff827b;
    assign coff[1535] = 64'h00001905ffff8278;
    assign coff[1536] = 64'h000018f9ffff8276;
    assign coff[1537] = 64'h000018ecffff8273;
    assign coff[1538] = 64'h000018e0ffff8271;
    assign coff[1539] = 64'h000018d4ffff826e;
    assign coff[1540] = 64'h000018c7ffff826c;
    assign coff[1541] = 64'h000018bbffff8269;
    assign coff[1542] = 64'h000018afffff8267;
    assign coff[1543] = 64'h000018a2ffff8265;
    assign coff[1544] = 64'h00001896ffff8262;
    assign coff[1545] = 64'h0000188affff8260;
    assign coff[1546] = 64'h0000187dffff825d;
    assign coff[1547] = 64'h00001871ffff825b;
    assign coff[1548] = 64'h00001865ffff8259;
    assign coff[1549] = 64'h00001858ffff8256;
    assign coff[1550] = 64'h0000184cffff8254;
    assign coff[1551] = 64'h00001840ffff8251;
    assign coff[1552] = 64'h00001833ffff824f;
    assign coff[1553] = 64'h00001827ffff824d;
    assign coff[1554] = 64'h0000181bffff824a;
    assign coff[1555] = 64'h0000180effff8248;
    assign coff[1556] = 64'h00001802ffff8246;
    assign coff[1557] = 64'h000017f6ffff8243;
    assign coff[1558] = 64'h000017e9ffff8241;
    assign coff[1559] = 64'h000017ddffff823e;
    assign coff[1560] = 64'h000017d1ffff823c;
    assign coff[1561] = 64'h000017c4ffff823a;
    assign coff[1562] = 64'h000017b8ffff8237;
    assign coff[1563] = 64'h000017acffff8235;
    assign coff[1564] = 64'h0000179fffff8233;
    assign coff[1565] = 64'h00001793ffff8231;
    assign coff[1566] = 64'h00001787ffff822e;
    assign coff[1567] = 64'h0000177affff822c;
    assign coff[1568] = 64'h0000176effff822a;
    assign coff[1569] = 64'h00001761ffff8227;
    assign coff[1570] = 64'h00001755ffff8225;
    assign coff[1571] = 64'h00001749ffff8223;
    assign coff[1572] = 64'h0000173cffff8220;
    assign coff[1573] = 64'h00001730ffff821e;
    assign coff[1574] = 64'h00001724ffff821c;
    assign coff[1575] = 64'h00001717ffff821a;
    assign coff[1576] = 64'h0000170bffff8217;
    assign coff[1577] = 64'h000016ffffff8215;
    assign coff[1578] = 64'h000016f2ffff8213;
    assign coff[1579] = 64'h000016e6ffff8211;
    assign coff[1580] = 64'h000016daffff820e;
    assign coff[1581] = 64'h000016cdffff820c;
    assign coff[1582] = 64'h000016c1ffff820a;
    assign coff[1583] = 64'h000016b4ffff8208;
    assign coff[1584] = 64'h000016a8ffff8205;
    assign coff[1585] = 64'h0000169cffff8203;
    assign coff[1586] = 64'h0000168fffff8201;
    assign coff[1587] = 64'h00001683ffff81ff;
    assign coff[1588] = 64'h00001677ffff81fd;
    assign coff[1589] = 64'h0000166affff81fa;
    assign coff[1590] = 64'h0000165effff81f8;
    assign coff[1591] = 64'h00001651ffff81f6;
    assign coff[1592] = 64'h00001645ffff81f4;
    assign coff[1593] = 64'h00001639ffff81f2;
    assign coff[1594] = 64'h0000162cffff81ef;
    assign coff[1595] = 64'h00001620ffff81ed;
    assign coff[1596] = 64'h00001614ffff81eb;
    assign coff[1597] = 64'h00001607ffff81e9;
    assign coff[1598] = 64'h000015fbffff81e7;
    assign coff[1599] = 64'h000015eeffff81e5;
    assign coff[1600] = 64'h000015e2ffff81e2;
    assign coff[1601] = 64'h000015d6ffff81e0;
    assign coff[1602] = 64'h000015c9ffff81de;
    assign coff[1603] = 64'h000015bdffff81dc;
    assign coff[1604] = 64'h000015b1ffff81da;
    assign coff[1605] = 64'h000015a4ffff81d8;
    assign coff[1606] = 64'h00001598ffff81d6;
    assign coff[1607] = 64'h0000158bffff81d3;
    assign coff[1608] = 64'h0000157fffff81d1;
    assign coff[1609] = 64'h00001573ffff81cf;
    assign coff[1610] = 64'h00001566ffff81cd;
    assign coff[1611] = 64'h0000155affff81cb;
    assign coff[1612] = 64'h0000154dffff81c9;
    assign coff[1613] = 64'h00001541ffff81c7;
    assign coff[1614] = 64'h00001535ffff81c5;
    assign coff[1615] = 64'h00001528ffff81c3;
    assign coff[1616] = 64'h0000151cffff81c1;
    assign coff[1617] = 64'h0000150fffff81bf;
    assign coff[1618] = 64'h00001503ffff81bd;
    assign coff[1619] = 64'h000014f7ffff81ba;
    assign coff[1620] = 64'h000014eaffff81b8;
    assign coff[1621] = 64'h000014deffff81b6;
    assign coff[1622] = 64'h000014d1ffff81b4;
    assign coff[1623] = 64'h000014c5ffff81b2;
    assign coff[1624] = 64'h000014b9ffff81b0;
    assign coff[1625] = 64'h000014acffff81ae;
    assign coff[1626] = 64'h000014a0ffff81ac;
    assign coff[1627] = 64'h00001493ffff81aa;
    assign coff[1628] = 64'h00001487ffff81a8;
    assign coff[1629] = 64'h0000147bffff81a6;
    assign coff[1630] = 64'h0000146effff81a4;
    assign coff[1631] = 64'h00001462ffff81a2;
    assign coff[1632] = 64'h00001455ffff81a0;
    assign coff[1633] = 64'h00001449ffff819e;
    assign coff[1634] = 64'h0000143dffff819c;
    assign coff[1635] = 64'h00001430ffff819a;
    assign coff[1636] = 64'h00001424ffff8198;
    assign coff[1637] = 64'h00001417ffff8196;
    assign coff[1638] = 64'h0000140bffff8194;
    assign coff[1639] = 64'h000013ffffff8192;
    assign coff[1640] = 64'h000013f2ffff8190;
    assign coff[1641] = 64'h000013e6ffff818e;
    assign coff[1642] = 64'h000013d9ffff818c;
    assign coff[1643] = 64'h000013cdffff818a;
    assign coff[1644] = 64'h000013c1ffff8188;
    assign coff[1645] = 64'h000013b4ffff8187;
    assign coff[1646] = 64'h000013a8ffff8185;
    assign coff[1647] = 64'h0000139bffff8183;
    assign coff[1648] = 64'h0000138fffff8181;
    assign coff[1649] = 64'h00001382ffff817f;
    assign coff[1650] = 64'h00001376ffff817d;
    assign coff[1651] = 64'h0000136affff817b;
    assign coff[1652] = 64'h0000135dffff8179;
    assign coff[1653] = 64'h00001351ffff8177;
    assign coff[1654] = 64'h00001344ffff8175;
    assign coff[1655] = 64'h00001338ffff8173;
    assign coff[1656] = 64'h0000132bffff8172;
    assign coff[1657] = 64'h0000131fffff8170;
    assign coff[1658] = 64'h00001313ffff816e;
    assign coff[1659] = 64'h00001306ffff816c;
    assign coff[1660] = 64'h000012faffff816a;
    assign coff[1661] = 64'h000012edffff8168;
    assign coff[1662] = 64'h000012e1ffff8166;
    assign coff[1663] = 64'h000012d4ffff8165;
    assign coff[1664] = 64'h000012c8ffff8163;
    assign coff[1665] = 64'h000012bcffff8161;
    assign coff[1666] = 64'h000012afffff815f;
    assign coff[1667] = 64'h000012a3ffff815d;
    assign coff[1668] = 64'h00001296ffff815b;
    assign coff[1669] = 64'h0000128affff815a;
    assign coff[1670] = 64'h0000127dffff8158;
    assign coff[1671] = 64'h00001271ffff8156;
    assign coff[1672] = 64'h00001265ffff8154;
    assign coff[1673] = 64'h00001258ffff8152;
    assign coff[1674] = 64'h0000124cffff8150;
    assign coff[1675] = 64'h0000123fffff814f;
    assign coff[1676] = 64'h00001233ffff814d;
    assign coff[1677] = 64'h00001226ffff814b;
    assign coff[1678] = 64'h0000121affff8149;
    assign coff[1679] = 64'h0000120effff8148;
    assign coff[1680] = 64'h00001201ffff8146;
    assign coff[1681] = 64'h000011f5ffff8144;
    assign coff[1682] = 64'h000011e8ffff8142;
    assign coff[1683] = 64'h000011dcffff8140;
    assign coff[1684] = 64'h000011cfffff813f;
    assign coff[1685] = 64'h000011c3ffff813d;
    assign coff[1686] = 64'h000011b6ffff813b;
    assign coff[1687] = 64'h000011aaffff813a;
    assign coff[1688] = 64'h0000119effff8138;
    assign coff[1689] = 64'h00001191ffff8136;
    assign coff[1690] = 64'h00001185ffff8134;
    assign coff[1691] = 64'h00001178ffff8133;
    assign coff[1692] = 64'h0000116cffff8131;
    assign coff[1693] = 64'h0000115fffff812f;
    assign coff[1694] = 64'h00001153ffff812d;
    assign coff[1695] = 64'h00001146ffff812c;
    assign coff[1696] = 64'h0000113affff812a;
    assign coff[1697] = 64'h0000112dffff8128;
    assign coff[1698] = 64'h00001121ffff8127;
    assign coff[1699] = 64'h00001115ffff8125;
    assign coff[1700] = 64'h00001108ffff8123;
    assign coff[1701] = 64'h000010fcffff8122;
    assign coff[1702] = 64'h000010efffff8120;
    assign coff[1703] = 64'h000010e3ffff811e;
    assign coff[1704] = 64'h000010d6ffff811d;
    assign coff[1705] = 64'h000010caffff811b;
    assign coff[1706] = 64'h000010bdffff8119;
    assign coff[1707] = 64'h000010b1ffff8118;
    assign coff[1708] = 64'h000010a4ffff8116;
    assign coff[1709] = 64'h00001098ffff8115;
    assign coff[1710] = 64'h0000108cffff8113;
    assign coff[1711] = 64'h0000107fffff8111;
    assign coff[1712] = 64'h00001073ffff8110;
    assign coff[1713] = 64'h00001066ffff810e;
    assign coff[1714] = 64'h0000105affff810c;
    assign coff[1715] = 64'h0000104dffff810b;
    assign coff[1716] = 64'h00001041ffff8109;
    assign coff[1717] = 64'h00001034ffff8108;
    assign coff[1718] = 64'h00001028ffff8106;
    assign coff[1719] = 64'h0000101bffff8104;
    assign coff[1720] = 64'h0000100fffff8103;
    assign coff[1721] = 64'h00001002ffff8101;
    assign coff[1722] = 64'h00000ff6ffff8100;
    assign coff[1723] = 64'h00000feaffff80fe;
    assign coff[1724] = 64'h00000fddffff80fd;
    assign coff[1725] = 64'h00000fd1ffff80fb;
    assign coff[1726] = 64'h00000fc4ffff80fa;
    assign coff[1727] = 64'h00000fb8ffff80f8;
    assign coff[1728] = 64'h00000fabffff80f6;
    assign coff[1729] = 64'h00000f9fffff80f5;
    assign coff[1730] = 64'h00000f92ffff80f3;
    assign coff[1731] = 64'h00000f86ffff80f2;
    assign coff[1732] = 64'h00000f79ffff80f0;
    assign coff[1733] = 64'h00000f6dffff80ef;
    assign coff[1734] = 64'h00000f60ffff80ed;
    assign coff[1735] = 64'h00000f54ffff80ec;
    assign coff[1736] = 64'h00000f47ffff80ea;
    assign coff[1737] = 64'h00000f3bffff80e9;
    assign coff[1738] = 64'h00000f2effff80e7;
    assign coff[1739] = 64'h00000f22ffff80e6;
    assign coff[1740] = 64'h00000f15ffff80e4;
    assign coff[1741] = 64'h00000f09ffff80e3;
    assign coff[1742] = 64'h00000efcffff80e1;
    assign coff[1743] = 64'h00000ef0ffff80e0;
    assign coff[1744] = 64'h00000ee4ffff80de;
    assign coff[1745] = 64'h00000ed7ffff80dd;
    assign coff[1746] = 64'h00000ecbffff80dc;
    assign coff[1747] = 64'h00000ebeffff80da;
    assign coff[1748] = 64'h00000eb2ffff80d9;
    assign coff[1749] = 64'h00000ea5ffff80d7;
    assign coff[1750] = 64'h00000e99ffff80d6;
    assign coff[1751] = 64'h00000e8cffff80d4;
    assign coff[1752] = 64'h00000e80ffff80d3;
    assign coff[1753] = 64'h00000e73ffff80d1;
    assign coff[1754] = 64'h00000e67ffff80d0;
    assign coff[1755] = 64'h00000e5affff80cf;
    assign coff[1756] = 64'h00000e4effff80cd;
    assign coff[1757] = 64'h00000e41ffff80cc;
    assign coff[1758] = 64'h00000e35ffff80ca;
    assign coff[1759] = 64'h00000e28ffff80c9;
    assign coff[1760] = 64'h00000e1cffff80c8;
    assign coff[1761] = 64'h00000e0fffff80c6;
    assign coff[1762] = 64'h00000e03ffff80c5;
    assign coff[1763] = 64'h00000df6ffff80c4;
    assign coff[1764] = 64'h00000deaffff80c2;
    assign coff[1765] = 64'h00000dddffff80c1;
    assign coff[1766] = 64'h00000dd1ffff80bf;
    assign coff[1767] = 64'h00000dc4ffff80be;
    assign coff[1768] = 64'h00000db8ffff80bd;
    assign coff[1769] = 64'h00000dabffff80bb;
    assign coff[1770] = 64'h00000d9fffff80ba;
    assign coff[1771] = 64'h00000d92ffff80b9;
    assign coff[1772] = 64'h00000d86ffff80b7;
    assign coff[1773] = 64'h00000d79ffff80b6;
    assign coff[1774] = 64'h00000d6dffff80b5;
    assign coff[1775] = 64'h00000d60ffff80b3;
    assign coff[1776] = 64'h00000d54ffff80b2;
    assign coff[1777] = 64'h00000d47ffff80b1;
    assign coff[1778] = 64'h00000d3bffff80b0;
    assign coff[1779] = 64'h00000d2effff80ae;
    assign coff[1780] = 64'h00000d22ffff80ad;
    assign coff[1781] = 64'h00000d15ffff80ac;
    assign coff[1782] = 64'h00000d09ffff80aa;
    assign coff[1783] = 64'h00000cfcffff80a9;
    assign coff[1784] = 64'h00000cf0ffff80a8;
    assign coff[1785] = 64'h00000ce3ffff80a7;
    assign coff[1786] = 64'h00000cd7ffff80a5;
    assign coff[1787] = 64'h00000ccaffff80a4;
    assign coff[1788] = 64'h00000cbeffff80a3;
    assign coff[1789] = 64'h00000cb1ffff80a2;
    assign coff[1790] = 64'h00000ca5ffff80a0;
    assign coff[1791] = 64'h00000c98ffff809f;
    assign coff[1792] = 64'h00000c8cffff809e;
    assign coff[1793] = 64'h00000c7fffff809d;
    assign coff[1794] = 64'h00000c73ffff809b;
    assign coff[1795] = 64'h00000c66ffff809a;
    assign coff[1796] = 64'h00000c5affff8099;
    assign coff[1797] = 64'h00000c4dffff8098;
    assign coff[1798] = 64'h00000c41ffff8096;
    assign coff[1799] = 64'h00000c34ffff8095;
    assign coff[1800] = 64'h00000c28ffff8094;
    assign coff[1801] = 64'h00000c1bffff8093;
    assign coff[1802] = 64'h00000c0fffff8092;
    assign coff[1803] = 64'h00000c02ffff8091;
    assign coff[1804] = 64'h00000bf6ffff808f;
    assign coff[1805] = 64'h00000be9ffff808e;
    assign coff[1806] = 64'h00000bddffff808d;
    assign coff[1807] = 64'h00000bd0ffff808c;
    assign coff[1808] = 64'h00000bc4ffff808b;
    assign coff[1809] = 64'h00000bb7ffff808a;
    assign coff[1810] = 64'h00000babffff8088;
    assign coff[1811] = 64'h00000b9effff8087;
    assign coff[1812] = 64'h00000b92ffff8086;
    assign coff[1813] = 64'h00000b85ffff8085;
    assign coff[1814] = 64'h00000b79ffff8084;
    assign coff[1815] = 64'h00000b6cffff8083;
    assign coff[1816] = 64'h00000b60ffff8082;
    assign coff[1817] = 64'h00000b53ffff8080;
    assign coff[1818] = 64'h00000b47ffff807f;
    assign coff[1819] = 64'h00000b3affff807e;
    assign coff[1820] = 64'h00000b2dffff807d;
    assign coff[1821] = 64'h00000b21ffff807c;
    assign coff[1822] = 64'h00000b14ffff807b;
    assign coff[1823] = 64'h00000b08ffff807a;
    assign coff[1824] = 64'h00000afbffff8079;
    assign coff[1825] = 64'h00000aefffff8078;
    assign coff[1826] = 64'h00000ae2ffff8077;
    assign coff[1827] = 64'h00000ad6ffff8076;
    assign coff[1828] = 64'h00000ac9ffff8075;
    assign coff[1829] = 64'h00000abdffff8073;
    assign coff[1830] = 64'h00000ab0ffff8072;
    assign coff[1831] = 64'h00000aa4ffff8071;
    assign coff[1832] = 64'h00000a97ffff8070;
    assign coff[1833] = 64'h00000a8bffff806f;
    assign coff[1834] = 64'h00000a7effff806e;
    assign coff[1835] = 64'h00000a72ffff806d;
    assign coff[1836] = 64'h00000a65ffff806c;
    assign coff[1837] = 64'h00000a59ffff806b;
    assign coff[1838] = 64'h00000a4cffff806a;
    assign coff[1839] = 64'h00000a40ffff8069;
    assign coff[1840] = 64'h00000a33ffff8068;
    assign coff[1841] = 64'h00000a27ffff8067;
    assign coff[1842] = 64'h00000a1affff8066;
    assign coff[1843] = 64'h00000a0dffff8065;
    assign coff[1844] = 64'h00000a01ffff8064;
    assign coff[1845] = 64'h000009f4ffff8063;
    assign coff[1846] = 64'h000009e8ffff8062;
    assign coff[1847] = 64'h000009dbffff8061;
    assign coff[1848] = 64'h000009cfffff8060;
    assign coff[1849] = 64'h000009c2ffff805f;
    assign coff[1850] = 64'h000009b6ffff805e;
    assign coff[1851] = 64'h000009a9ffff805d;
    assign coff[1852] = 64'h0000099dffff805d;
    assign coff[1853] = 64'h00000990ffff805c;
    assign coff[1854] = 64'h00000984ffff805b;
    assign coff[1855] = 64'h00000977ffff805a;
    assign coff[1856] = 64'h0000096bffff8059;
    assign coff[1857] = 64'h0000095effff8058;
    assign coff[1858] = 64'h00000951ffff8057;
    assign coff[1859] = 64'h00000945ffff8056;
    assign coff[1860] = 64'h00000938ffff8055;
    assign coff[1861] = 64'h0000092cffff8054;
    assign coff[1862] = 64'h0000091fffff8053;
    assign coff[1863] = 64'h00000913ffff8052;
    assign coff[1864] = 64'h00000906ffff8052;
    assign coff[1865] = 64'h000008faffff8051;
    assign coff[1866] = 64'h000008edffff8050;
    assign coff[1867] = 64'h000008e1ffff804f;
    assign coff[1868] = 64'h000008d4ffff804e;
    assign coff[1869] = 64'h000008c8ffff804d;
    assign coff[1870] = 64'h000008bbffff804c;
    assign coff[1871] = 64'h000008afffff804b;
    assign coff[1872] = 64'h000008a2ffff804b;
    assign coff[1873] = 64'h00000895ffff804a;
    assign coff[1874] = 64'h00000889ffff8049;
    assign coff[1875] = 64'h0000087cffff8048;
    assign coff[1876] = 64'h00000870ffff8047;
    assign coff[1877] = 64'h00000863ffff8046;
    assign coff[1878] = 64'h00000857ffff8046;
    assign coff[1879] = 64'h0000084affff8045;
    assign coff[1880] = 64'h0000083effff8044;
    assign coff[1881] = 64'h00000831ffff8043;
    assign coff[1882] = 64'h00000825ffff8042;
    assign coff[1883] = 64'h00000818ffff8042;
    assign coff[1884] = 64'h0000080cffff8041;
    assign coff[1885] = 64'h000007ffffff8040;
    assign coff[1886] = 64'h000007f2ffff803f;
    assign coff[1887] = 64'h000007e6ffff803e;
    assign coff[1888] = 64'h000007d9ffff803e;
    assign coff[1889] = 64'h000007cdffff803d;
    assign coff[1890] = 64'h000007c0ffff803c;
    assign coff[1891] = 64'h000007b4ffff803b;
    assign coff[1892] = 64'h000007a7ffff803b;
    assign coff[1893] = 64'h0000079bffff803a;
    assign coff[1894] = 64'h0000078effff8039;
    assign coff[1895] = 64'h00000782ffff8038;
    assign coff[1896] = 64'h00000775ffff8038;
    assign coff[1897] = 64'h00000768ffff8037;
    assign coff[1898] = 64'h0000075cffff8036;
    assign coff[1899] = 64'h0000074fffff8035;
    assign coff[1900] = 64'h00000743ffff8035;
    assign coff[1901] = 64'h00000736ffff8034;
    assign coff[1902] = 64'h0000072affff8033;
    assign coff[1903] = 64'h0000071dffff8033;
    assign coff[1904] = 64'h00000711ffff8032;
    assign coff[1905] = 64'h00000704ffff8031;
    assign coff[1906] = 64'h000006f8ffff8031;
    assign coff[1907] = 64'h000006ebffff8030;
    assign coff[1908] = 64'h000006deffff802f;
    assign coff[1909] = 64'h000006d2ffff802f;
    assign coff[1910] = 64'h000006c5ffff802e;
    assign coff[1911] = 64'h000006b9ffff802d;
    assign coff[1912] = 64'h000006acffff802d;
    assign coff[1913] = 64'h000006a0ffff802c;
    assign coff[1914] = 64'h00000693ffff802b;
    assign coff[1915] = 64'h00000687ffff802b;
    assign coff[1916] = 64'h0000067affff802a;
    assign coff[1917] = 64'h0000066effff8029;
    assign coff[1918] = 64'h00000661ffff8029;
    assign coff[1919] = 64'h00000654ffff8028;
    assign coff[1920] = 64'h00000648ffff8027;
    assign coff[1921] = 64'h0000063bffff8027;
    assign coff[1922] = 64'h0000062fffff8026;
    assign coff[1923] = 64'h00000622ffff8026;
    assign coff[1924] = 64'h00000616ffff8025;
    assign coff[1925] = 64'h00000609ffff8024;
    assign coff[1926] = 64'h000005fdffff8024;
    assign coff[1927] = 64'h000005f0ffff8023;
    assign coff[1928] = 64'h000005e3ffff8023;
    assign coff[1929] = 64'h000005d7ffff8022;
    assign coff[1930] = 64'h000005caffff8022;
    assign coff[1931] = 64'h000005beffff8021;
    assign coff[1932] = 64'h000005b1ffff8020;
    assign coff[1933] = 64'h000005a5ffff8020;
    assign coff[1934] = 64'h00000598ffff801f;
    assign coff[1935] = 64'h0000058cffff801f;
    assign coff[1936] = 64'h0000057fffff801e;
    assign coff[1937] = 64'h00000572ffff801e;
    assign coff[1938] = 64'h00000566ffff801d;
    assign coff[1939] = 64'h00000559ffff801d;
    assign coff[1940] = 64'h0000054dffff801c;
    assign coff[1941] = 64'h00000540ffff801c;
    assign coff[1942] = 64'h00000534ffff801b;
    assign coff[1943] = 64'h00000527ffff801b;
    assign coff[1944] = 64'h0000051bffff801a;
    assign coff[1945] = 64'h0000050effff801a;
    assign coff[1946] = 64'h00000501ffff8019;
    assign coff[1947] = 64'h000004f5ffff8019;
    assign coff[1948] = 64'h000004e8ffff8018;
    assign coff[1949] = 64'h000004dcffff8018;
    assign coff[1950] = 64'h000004cfffff8017;
    assign coff[1951] = 64'h000004c3ffff8017;
    assign coff[1952] = 64'h000004b6ffff8016;
    assign coff[1953] = 64'h000004aaffff8016;
    assign coff[1954] = 64'h0000049dffff8015;
    assign coff[1955] = 64'h00000490ffff8015;
    assign coff[1956] = 64'h00000484ffff8014;
    assign coff[1957] = 64'h00000477ffff8014;
    assign coff[1958] = 64'h0000046bffff8014;
    assign coff[1959] = 64'h0000045effff8013;
    assign coff[1960] = 64'h00000452ffff8013;
    assign coff[1961] = 64'h00000445ffff8012;
    assign coff[1962] = 64'h00000439ffff8012;
    assign coff[1963] = 64'h0000042cffff8011;
    assign coff[1964] = 64'h0000041fffff8011;
    assign coff[1965] = 64'h00000413ffff8011;
    assign coff[1966] = 64'h00000406ffff8010;
    assign coff[1967] = 64'h000003faffff8010;
    assign coff[1968] = 64'h000003edffff800f;
    assign coff[1969] = 64'h000003e1ffff800f;
    assign coff[1970] = 64'h000003d4ffff800f;
    assign coff[1971] = 64'h000003c7ffff800e;
    assign coff[1972] = 64'h000003bbffff800e;
    assign coff[1973] = 64'h000003aeffff800e;
    assign coff[1974] = 64'h000003a2ffff800d;
    assign coff[1975] = 64'h00000395ffff800d;
    assign coff[1976] = 64'h00000389ffff800c;
    assign coff[1977] = 64'h0000037cffff800c;
    assign coff[1978] = 64'h00000370ffff800c;
    assign coff[1979] = 64'h00000363ffff800b;
    assign coff[1980] = 64'h00000356ffff800b;
    assign coff[1981] = 64'h0000034affff800b;
    assign coff[1982] = 64'h0000033dffff800a;
    assign coff[1983] = 64'h00000331ffff800a;
    assign coff[1984] = 64'h00000324ffff800a;
    assign coff[1985] = 64'h00000318ffff800a;
    assign coff[1986] = 64'h0000030bffff8009;
    assign coff[1987] = 64'h000002feffff8009;
    assign coff[1988] = 64'h000002f2ffff8009;
    assign coff[1989] = 64'h000002e5ffff8008;
    assign coff[1990] = 64'h000002d9ffff8008;
    assign coff[1991] = 64'h000002ccffff8008;
    assign coff[1992] = 64'h000002c0ffff8008;
    assign coff[1993] = 64'h000002b3ffff8007;
    assign coff[1994] = 64'h000002a7ffff8007;
    assign coff[1995] = 64'h0000029affff8007;
    assign coff[1996] = 64'h0000028dffff8007;
    assign coff[1997] = 64'h00000281ffff8006;
    assign coff[1998] = 64'h00000274ffff8006;
    assign coff[1999] = 64'h00000268ffff8006;
    assign coff[2000] = 64'h0000025bffff8006;
    assign coff[2001] = 64'h0000024fffff8005;
    assign coff[2002] = 64'h00000242ffff8005;
    assign coff[2003] = 64'h00000235ffff8005;
    assign coff[2004] = 64'h00000229ffff8005;
    assign coff[2005] = 64'h0000021cffff8004;
    assign coff[2006] = 64'h00000210ffff8004;
    assign coff[2007] = 64'h00000203ffff8004;
    assign coff[2008] = 64'h000001f7ffff8004;
    assign coff[2009] = 64'h000001eaffff8004;
    assign coff[2010] = 64'h000001deffff8003;
    assign coff[2011] = 64'h000001d1ffff8003;
    assign coff[2012] = 64'h000001c4ffff8003;
    assign coff[2013] = 64'h000001b8ffff8003;
    assign coff[2014] = 64'h000001abffff8003;
    assign coff[2015] = 64'h0000019fffff8003;
    assign coff[2016] = 64'h00000192ffff8002;
    assign coff[2017] = 64'h00000186ffff8002;
    assign coff[2018] = 64'h00000179ffff8002;
    assign coff[2019] = 64'h0000016cffff8002;
    assign coff[2020] = 64'h00000160ffff8002;
    assign coff[2021] = 64'h00000153ffff8002;
    assign coff[2022] = 64'h00000147ffff8002;
    assign coff[2023] = 64'h0000013affff8002;
    assign coff[2024] = 64'h0000012effff8001;
    assign coff[2025] = 64'h00000121ffff8001;
    assign coff[2026] = 64'h00000114ffff8001;
    assign coff[2027] = 64'h00000108ffff8001;
    assign coff[2028] = 64'h000000fbffff8001;
    assign coff[2029] = 64'h000000efffff8001;
    assign coff[2030] = 64'h000000e2ffff8001;
    assign coff[2031] = 64'h000000d6ffff8001;
    assign coff[2032] = 64'h000000c9ffff8001;
    assign coff[2033] = 64'h000000bcffff8001;
    assign coff[2034] = 64'h000000b0ffff8001;
    assign coff[2035] = 64'h000000a3ffff8001;
    assign coff[2036] = 64'h00000097ffff8001;
    assign coff[2037] = 64'h0000008affff8001;
    assign coff[2038] = 64'h0000007effff8001;
    assign coff[2039] = 64'h00000071ffff8001;
    assign coff[2040] = 64'h00000065ffff8001;
    assign coff[2041] = 64'h00000058ffff8001;
    assign coff[2042] = 64'h0000004bffff8001;
    assign coff[2043] = 64'h0000003fffff8001;
    assign coff[2044] = 64'h00000032ffff8001;
    assign coff[2045] = 64'h00000026ffff8001;
    assign coff[2046] = 64'h00000019ffff8001;
    assign coff[2047] = 64'h0000000dffff8001;




    always_ff @(posedge clk, negedge rst_n) begin
        if(~rst_n) begin
            data_o_col1 <= 'b0;
            data_o_col2 <= 'b0;
        end else begin
            if ((addr_col1 == 'd0 || addr_col1 == 'd1024) && (valid == 1)) begin
                data_o_col1 <= coff[addr_col1];
                data_o_col2 <= 'b0;
            end else if(valid == 1) begin
                data_o_col1 <= coff[addr_col1];
                data_o_col2 <= coff[addr_col2];
            end else begin
                data_o_col1 <= 'b0;
                data_o_col2 <= 'b0;
            end       
        end
    end


endmodule