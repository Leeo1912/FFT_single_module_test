// `timescale 1ns/1ps
module rom_3_rfft_data64
(
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic                     valid,
    input  logic [10:0]              addr_col1,
    input  logic [10:0]              addr_col2,
    output logic [63:0]              data_o_col1,
    output logic [63:0]              data_o_col2
);

    logic [63:0] coff[2047:0];

    assign coff[0   ] = 64'h00000000ffff8001;
    assign coff[1   ] = 64'hfffffff3ffff8001;
    assign coff[2   ] = 64'hffffffe7ffff8001;
    assign coff[3   ] = 64'hffffffdaffff8001;
    assign coff[4   ] = 64'hffffffceffff8001;
    assign coff[5   ] = 64'hffffffc1ffff8001;
    assign coff[6   ] = 64'hffffffb5ffff8001;
    assign coff[7   ] = 64'hffffffa8ffff8001;
    assign coff[8   ] = 64'hffffff9bffff8001;
    assign coff[9   ] = 64'hffffff8fffff8001;
    assign coff[10  ] = 64'hffffff82ffff8001;
    assign coff[11  ] = 64'hffffff76ffff8001;
    assign coff[12  ] = 64'hffffff69ffff8001;
    assign coff[13  ] = 64'hffffff5dffff8001;
    assign coff[14  ] = 64'hffffff50ffff8001;
    assign coff[15  ] = 64'hffffff44ffff8001;
    assign coff[16  ] = 64'hffffff37ffff8001;
    assign coff[17  ] = 64'hffffff2affff8001;
    assign coff[18  ] = 64'hffffff1effff8001;
    assign coff[19  ] = 64'hffffff11ffff8001;
    assign coff[20  ] = 64'hffffff05ffff8001;
    assign coff[21  ] = 64'hfffffef8ffff8001;
    assign coff[22  ] = 64'hfffffeecffff8001;
    assign coff[23  ] = 64'hfffffedfffff8001;
    assign coff[24  ] = 64'hfffffed2ffff8001;
    assign coff[25  ] = 64'hfffffec6ffff8002;
    assign coff[26  ] = 64'hfffffeb9ffff8002;
    assign coff[27  ] = 64'hfffffeadffff8002;
    assign coff[28  ] = 64'hfffffea0ffff8002;
    assign coff[29  ] = 64'hfffffe94ffff8002;
    assign coff[30  ] = 64'hfffffe87ffff8002;
    assign coff[31  ] = 64'hfffffe7affff8002;
    assign coff[32  ] = 64'hfffffe6effff8002;
    assign coff[33  ] = 64'hfffffe61ffff8003;
    assign coff[34  ] = 64'hfffffe55ffff8003;
    assign coff[35  ] = 64'hfffffe48ffff8003;
    assign coff[36  ] = 64'hfffffe3cffff8003;
    assign coff[37  ] = 64'hfffffe2fffff8003;
    assign coff[38  ] = 64'hfffffe22ffff8003;
    assign coff[39  ] = 64'hfffffe16ffff8004;
    assign coff[40  ] = 64'hfffffe09ffff8004;
    assign coff[41  ] = 64'hfffffdfdffff8004;
    assign coff[42  ] = 64'hfffffdf0ffff8004;
    assign coff[43  ] = 64'hfffffde4ffff8004;
    assign coff[44  ] = 64'hfffffdd7ffff8005;
    assign coff[45  ] = 64'hfffffdcbffff8005;
    assign coff[46  ] = 64'hfffffdbeffff8005;
    assign coff[47  ] = 64'hfffffdb1ffff8005;
    assign coff[48  ] = 64'hfffffda5ffff8006;
    assign coff[49  ] = 64'hfffffd98ffff8006;
    assign coff[50  ] = 64'hfffffd8cffff8006;
    assign coff[51  ] = 64'hfffffd7fffff8006;
    assign coff[52  ] = 64'hfffffd73ffff8007;
    assign coff[53  ] = 64'hfffffd66ffff8007;
    assign coff[54  ] = 64'hfffffd59ffff8007;
    assign coff[55  ] = 64'hfffffd4dffff8007;
    assign coff[56  ] = 64'hfffffd40ffff8008;
    assign coff[57  ] = 64'hfffffd34ffff8008;
    assign coff[58  ] = 64'hfffffd27ffff8008;
    assign coff[59  ] = 64'hfffffd1bffff8008;
    assign coff[60  ] = 64'hfffffd0effff8009;
    assign coff[61  ] = 64'hfffffd02ffff8009;
    assign coff[62  ] = 64'hfffffcf5ffff8009;
    assign coff[63  ] = 64'hfffffce8ffff800a;
    assign coff[64  ] = 64'hfffffcdcffff800a;
    assign coff[65  ] = 64'hfffffccfffff800a;
    assign coff[66  ] = 64'hfffffcc3ffff800a;
    assign coff[67  ] = 64'hfffffcb6ffff800b;
    assign coff[68  ] = 64'hfffffcaaffff800b;
    assign coff[69  ] = 64'hfffffc9dffff800b;
    assign coff[70  ] = 64'hfffffc90ffff800c;
    assign coff[71  ] = 64'hfffffc84ffff800c;
    assign coff[72  ] = 64'hfffffc77ffff800c;
    assign coff[73  ] = 64'hfffffc6bffff800d;
    assign coff[74  ] = 64'hfffffc5effff800d;
    assign coff[75  ] = 64'hfffffc52ffff800e;
    assign coff[76  ] = 64'hfffffc45ffff800e;
    assign coff[77  ] = 64'hfffffc39ffff800e;
    assign coff[78  ] = 64'hfffffc2cffff800f;
    assign coff[79  ] = 64'hfffffc1fffff800f;
    assign coff[80  ] = 64'hfffffc13ffff800f;
    assign coff[81  ] = 64'hfffffc06ffff8010;
    assign coff[82  ] = 64'hfffffbfaffff8010;
    assign coff[83  ] = 64'hfffffbedffff8011;
    assign coff[84  ] = 64'hfffffbe1ffff8011;
    assign coff[85  ] = 64'hfffffbd4ffff8011;
    assign coff[86  ] = 64'hfffffbc7ffff8012;
    assign coff[87  ] = 64'hfffffbbbffff8012;
    assign coff[88  ] = 64'hfffffbaeffff8013;
    assign coff[89  ] = 64'hfffffba2ffff8013;
    assign coff[90  ] = 64'hfffffb95ffff8014;
    assign coff[91  ] = 64'hfffffb89ffff8014;
    assign coff[92  ] = 64'hfffffb7cffff8014;
    assign coff[93  ] = 64'hfffffb70ffff8015;
    assign coff[94  ] = 64'hfffffb63ffff8015;
    assign coff[95  ] = 64'hfffffb56ffff8016;
    assign coff[96  ] = 64'hfffffb4affff8016;
    assign coff[97  ] = 64'hfffffb3dffff8017;
    assign coff[98  ] = 64'hfffffb31ffff8017;
    assign coff[99  ] = 64'hfffffb24ffff8018;
    assign coff[100 ] = 64'hfffffb18ffff8018;
    assign coff[101 ] = 64'hfffffb0bffff8019;
    assign coff[102 ] = 64'hfffffaffffff8019;
    assign coff[103 ] = 64'hfffffaf2ffff801a;
    assign coff[104 ] = 64'hfffffae5ffff801a;
    assign coff[105 ] = 64'hfffffad9ffff801b;
    assign coff[106 ] = 64'hfffffaccffff801b;
    assign coff[107 ] = 64'hfffffac0ffff801c;
    assign coff[108 ] = 64'hfffffab3ffff801c;
    assign coff[109 ] = 64'hfffffaa7ffff801d;
    assign coff[110 ] = 64'hfffffa9affff801d;
    assign coff[111 ] = 64'hfffffa8effff801e;
    assign coff[112 ] = 64'hfffffa81ffff801e;
    assign coff[113 ] = 64'hfffffa74ffff801f;
    assign coff[114 ] = 64'hfffffa68ffff801f;
    assign coff[115 ] = 64'hfffffa5bffff8020;
    assign coff[116 ] = 64'hfffffa4fffff8020;
    assign coff[117 ] = 64'hfffffa42ffff8021;
    assign coff[118 ] = 64'hfffffa36ffff8022;
    assign coff[119 ] = 64'hfffffa29ffff8022;
    assign coff[120 ] = 64'hfffffa1dffff8023;
    assign coff[121 ] = 64'hfffffa10ffff8023;
    assign coff[122 ] = 64'hfffffa03ffff8024;
    assign coff[123 ] = 64'hfffff9f7ffff8024;
    assign coff[124 ] = 64'hfffff9eaffff8025;
    assign coff[125 ] = 64'hfffff9deffff8026;
    assign coff[126 ] = 64'hfffff9d1ffff8026;
    assign coff[127 ] = 64'hfffff9c5ffff8027;
    assign coff[128 ] = 64'hfffff9b8ffff8027;
    assign coff[129 ] = 64'hfffff9acffff8028;
    assign coff[130 ] = 64'hfffff99fffff8029;
    assign coff[131 ] = 64'hfffff992ffff8029;
    assign coff[132 ] = 64'hfffff986ffff802a;
    assign coff[133 ] = 64'hfffff979ffff802b;
    assign coff[134 ] = 64'hfffff96dffff802b;
    assign coff[135 ] = 64'hfffff960ffff802c;
    assign coff[136 ] = 64'hfffff954ffff802d;
    assign coff[137 ] = 64'hfffff947ffff802d;
    assign coff[138 ] = 64'hfffff93bffff802e;
    assign coff[139 ] = 64'hfffff92effff802f;
    assign coff[140 ] = 64'hfffff922ffff802f;
    assign coff[141 ] = 64'hfffff915ffff8030;
    assign coff[142 ] = 64'hfffff908ffff8031;
    assign coff[143 ] = 64'hfffff8fcffff8031;
    assign coff[144 ] = 64'hfffff8efffff8032;
    assign coff[145 ] = 64'hfffff8e3ffff8033;
    assign coff[146 ] = 64'hfffff8d6ffff8033;
    assign coff[147 ] = 64'hfffff8caffff8034;
    assign coff[148 ] = 64'hfffff8bdffff8035;
    assign coff[149 ] = 64'hfffff8b1ffff8035;
    assign coff[150 ] = 64'hfffff8a4ffff8036;
    assign coff[151 ] = 64'hfffff898ffff8037;
    assign coff[152 ] = 64'hfffff88bffff8038;
    assign coff[153 ] = 64'hfffff87effff8038;
    assign coff[154 ] = 64'hfffff872ffff8039;
    assign coff[155 ] = 64'hfffff865ffff803a;
    assign coff[156 ] = 64'hfffff859ffff803b;
    assign coff[157 ] = 64'hfffff84cffff803b;
    assign coff[158 ] = 64'hfffff840ffff803c;
    assign coff[159 ] = 64'hfffff833ffff803d;
    assign coff[160 ] = 64'hfffff827ffff803e;
    assign coff[161 ] = 64'hfffff81affff803e;
    assign coff[162 ] = 64'hfffff80effff803f;
    assign coff[163 ] = 64'hfffff801ffff8040;
    assign coff[164 ] = 64'hfffff7f4ffff8041;
    assign coff[165 ] = 64'hfffff7e8ffff8042;
    assign coff[166 ] = 64'hfffff7dbffff8042;
    assign coff[167 ] = 64'hfffff7cfffff8043;
    assign coff[168 ] = 64'hfffff7c2ffff8044;
    assign coff[169 ] = 64'hfffff7b6ffff8045;
    assign coff[170 ] = 64'hfffff7a9ffff8046;
    assign coff[171 ] = 64'hfffff79dffff8046;
    assign coff[172 ] = 64'hfffff790ffff8047;
    assign coff[173 ] = 64'hfffff784ffff8048;
    assign coff[174 ] = 64'hfffff777ffff8049;
    assign coff[175 ] = 64'hfffff76bffff804a;
    assign coff[176 ] = 64'hfffff75effff804b;
    assign coff[177 ] = 64'hfffff751ffff804b;
    assign coff[178 ] = 64'hfffff745ffff804c;
    assign coff[179 ] = 64'hfffff738ffff804d;
    assign coff[180 ] = 64'hfffff72cffff804e;
    assign coff[181 ] = 64'hfffff71fffff804f;
    assign coff[182 ] = 64'hfffff713ffff8050;
    assign coff[183 ] = 64'hfffff706ffff8051;
    assign coff[184 ] = 64'hfffff6faffff8052;
    assign coff[185 ] = 64'hfffff6edffff8052;
    assign coff[186 ] = 64'hfffff6e1ffff8053;
    assign coff[187 ] = 64'hfffff6d4ffff8054;
    assign coff[188 ] = 64'hfffff6c8ffff8055;
    assign coff[189 ] = 64'hfffff6bbffff8056;
    assign coff[190 ] = 64'hfffff6afffff8057;
    assign coff[191 ] = 64'hfffff6a2ffff8058;
    assign coff[192 ] = 64'hfffff695ffff8059;
    assign coff[193 ] = 64'hfffff689ffff805a;
    assign coff[194 ] = 64'hfffff67cffff805b;
    assign coff[195 ] = 64'hfffff670ffff805c;
    assign coff[196 ] = 64'hfffff663ffff805d;
    assign coff[197 ] = 64'hfffff657ffff805d;
    assign coff[198 ] = 64'hfffff64affff805e;
    assign coff[199 ] = 64'hfffff63effff805f;
    assign coff[200 ] = 64'hfffff631ffff8060;
    assign coff[201 ] = 64'hfffff625ffff8061;
    assign coff[202 ] = 64'hfffff618ffff8062;
    assign coff[203 ] = 64'hfffff60cffff8063;
    assign coff[204 ] = 64'hfffff5ffffff8064;
    assign coff[205 ] = 64'hfffff5f3ffff8065;
    assign coff[206 ] = 64'hfffff5e6ffff8066;
    assign coff[207 ] = 64'hfffff5d9ffff8067;
    assign coff[208 ] = 64'hfffff5cdffff8068;
    assign coff[209 ] = 64'hfffff5c0ffff8069;
    assign coff[210 ] = 64'hfffff5b4ffff806a;
    assign coff[211 ] = 64'hfffff5a7ffff806b;
    assign coff[212 ] = 64'hfffff59bffff806c;
    assign coff[213 ] = 64'hfffff58effff806d;
    assign coff[214 ] = 64'hfffff582ffff806e;
    assign coff[215 ] = 64'hfffff575ffff806f;
    assign coff[216 ] = 64'hfffff569ffff8070;
    assign coff[217 ] = 64'hfffff55cffff8071;
    assign coff[218 ] = 64'hfffff550ffff8072;
    assign coff[219 ] = 64'hfffff543ffff8073;
    assign coff[220 ] = 64'hfffff537ffff8075;
    assign coff[221 ] = 64'hfffff52affff8076;
    assign coff[222 ] = 64'hfffff51effff8077;
    assign coff[223 ] = 64'hfffff511ffff8078;
    assign coff[224 ] = 64'hfffff505ffff8079;
    assign coff[225 ] = 64'hfffff4f8ffff807a;
    assign coff[226 ] = 64'hfffff4ecffff807b;
    assign coff[227 ] = 64'hfffff4dfffff807c;
    assign coff[228 ] = 64'hfffff4d3ffff807d;
    assign coff[229 ] = 64'hfffff4c6ffff807e;
    assign coff[230 ] = 64'hfffff4b9ffff807f;
    assign coff[231 ] = 64'hfffff4adffff8080;
    assign coff[232 ] = 64'hfffff4a0ffff8082;
    assign coff[233 ] = 64'hfffff494ffff8083;
    assign coff[234 ] = 64'hfffff487ffff8084;
    assign coff[235 ] = 64'hfffff47bffff8085;
    assign coff[236 ] = 64'hfffff46effff8086;
    assign coff[237 ] = 64'hfffff462ffff8087;
    assign coff[238 ] = 64'hfffff455ffff8088;
    assign coff[239 ] = 64'hfffff449ffff808a;
    assign coff[240 ] = 64'hfffff43cffff808b;
    assign coff[241 ] = 64'hfffff430ffff808c;
    assign coff[242 ] = 64'hfffff423ffff808d;
    assign coff[243 ] = 64'hfffff417ffff808e;
    assign coff[244 ] = 64'hfffff40affff808f;
    assign coff[245 ] = 64'hfffff3feffff8091;
    assign coff[246 ] = 64'hfffff3f1ffff8092;
    assign coff[247 ] = 64'hfffff3e5ffff8093;
    assign coff[248 ] = 64'hfffff3d8ffff8094;
    assign coff[249 ] = 64'hfffff3ccffff8095;
    assign coff[250 ] = 64'hfffff3bfffff8096;
    assign coff[251 ] = 64'hfffff3b3ffff8098;
    assign coff[252 ] = 64'hfffff3a6ffff8099;
    assign coff[253 ] = 64'hfffff39affff809a;
    assign coff[254 ] = 64'hfffff38dffff809b;
    assign coff[255 ] = 64'hfffff381ffff809d;
    assign coff[256 ] = 64'hfffff374ffff809e;
    assign coff[257 ] = 64'hfffff368ffff809f;
    assign coff[258 ] = 64'hfffff35bffff80a0;
    assign coff[259 ] = 64'hfffff34fffff80a2;
    assign coff[260 ] = 64'hfffff342ffff80a3;
    assign coff[261 ] = 64'hfffff336ffff80a4;
    assign coff[262 ] = 64'hfffff329ffff80a5;
    assign coff[263 ] = 64'hfffff31dffff80a7;
    assign coff[264 ] = 64'hfffff310ffff80a8;
    assign coff[265 ] = 64'hfffff304ffff80a9;
    assign coff[266 ] = 64'hfffff2f7ffff80aa;
    assign coff[267 ] = 64'hfffff2ebffff80ac;
    assign coff[268 ] = 64'hfffff2deffff80ad;
    assign coff[269 ] = 64'hfffff2d2ffff80ae;
    assign coff[270 ] = 64'hfffff2c5ffff80b0;
    assign coff[271 ] = 64'hfffff2b9ffff80b1;
    assign coff[272 ] = 64'hfffff2acffff80b2;
    assign coff[273 ] = 64'hfffff2a0ffff80b3;
    assign coff[274 ] = 64'hfffff293ffff80b5;
    assign coff[275 ] = 64'hfffff287ffff80b6;
    assign coff[276 ] = 64'hfffff27affff80b7;
    assign coff[277 ] = 64'hfffff26effff80b9;
    assign coff[278 ] = 64'hfffff261ffff80ba;
    assign coff[279 ] = 64'hfffff255ffff80bb;
    assign coff[280 ] = 64'hfffff248ffff80bd;
    assign coff[281 ] = 64'hfffff23cffff80be;
    assign coff[282 ] = 64'hfffff22fffff80bf;
    assign coff[283 ] = 64'hfffff223ffff80c1;
    assign coff[284 ] = 64'hfffff216ffff80c2;
    assign coff[285 ] = 64'hfffff20affff80c4;
    assign coff[286 ] = 64'hfffff1fdffff80c5;
    assign coff[287 ] = 64'hfffff1f1ffff80c6;
    assign coff[288 ] = 64'hfffff1e4ffff80c8;
    assign coff[289 ] = 64'hfffff1d8ffff80c9;
    assign coff[290 ] = 64'hfffff1cbffff80ca;
    assign coff[291 ] = 64'hfffff1bfffff80cc;
    assign coff[292 ] = 64'hfffff1b2ffff80cd;
    assign coff[293 ] = 64'hfffff1a6ffff80cf;
    assign coff[294 ] = 64'hfffff199ffff80d0;
    assign coff[295 ] = 64'hfffff18dffff80d1;
    assign coff[296 ] = 64'hfffff180ffff80d3;
    assign coff[297 ] = 64'hfffff174ffff80d4;
    assign coff[298 ] = 64'hfffff167ffff80d6;
    assign coff[299 ] = 64'hfffff15bffff80d7;
    assign coff[300 ] = 64'hfffff14effff80d9;
    assign coff[301 ] = 64'hfffff142ffff80da;
    assign coff[302 ] = 64'hfffff135ffff80dc;
    assign coff[303 ] = 64'hfffff129ffff80dd;
    assign coff[304 ] = 64'hfffff11cffff80de;
    assign coff[305 ] = 64'hfffff110ffff80e0;
    assign coff[306 ] = 64'hfffff104ffff80e1;
    assign coff[307 ] = 64'hfffff0f7ffff80e3;
    assign coff[308 ] = 64'hfffff0ebffff80e4;
    assign coff[309 ] = 64'hfffff0deffff80e6;
    assign coff[310 ] = 64'hfffff0d2ffff80e7;
    assign coff[311 ] = 64'hfffff0c5ffff80e9;
    assign coff[312 ] = 64'hfffff0b9ffff80ea;
    assign coff[313 ] = 64'hfffff0acffff80ec;
    assign coff[314 ] = 64'hfffff0a0ffff80ed;
    assign coff[315 ] = 64'hfffff093ffff80ef;
    assign coff[316 ] = 64'hfffff087ffff80f0;
    assign coff[317 ] = 64'hfffff07affff80f2;
    assign coff[318 ] = 64'hfffff06effff80f3;
    assign coff[319 ] = 64'hfffff061ffff80f5;
    assign coff[320 ] = 64'hfffff055ffff80f6;
    assign coff[321 ] = 64'hfffff048ffff80f8;
    assign coff[322 ] = 64'hfffff03cffff80fa;
    assign coff[323 ] = 64'hfffff02fffff80fb;
    assign coff[324 ] = 64'hfffff023ffff80fd;
    assign coff[325 ] = 64'hfffff016ffff80fe;
    assign coff[326 ] = 64'hfffff00affff8100;
    assign coff[327 ] = 64'hffffeffeffff8101;
    assign coff[328 ] = 64'hffffeff1ffff8103;
    assign coff[329 ] = 64'hffffefe5ffff8104;
    assign coff[330 ] = 64'hffffefd8ffff8106;
    assign coff[331 ] = 64'hffffefccffff8108;
    assign coff[332 ] = 64'hffffefbfffff8109;
    assign coff[333 ] = 64'hffffefb3ffff810b;
    assign coff[334 ] = 64'hffffefa6ffff810c;
    assign coff[335 ] = 64'hffffef9affff810e;
    assign coff[336 ] = 64'hffffef8dffff8110;
    assign coff[337 ] = 64'hffffef81ffff8111;
    assign coff[338 ] = 64'hffffef74ffff8113;
    assign coff[339 ] = 64'hffffef68ffff8115;
    assign coff[340 ] = 64'hffffef5cffff8116;
    assign coff[341 ] = 64'hffffef4fffff8118;
    assign coff[342 ] = 64'hffffef43ffff8119;
    assign coff[343 ] = 64'hffffef36ffff811b;
    assign coff[344 ] = 64'hffffef2affff811d;
    assign coff[345 ] = 64'hffffef1dffff811e;
    assign coff[346 ] = 64'hffffef11ffff8120;
    assign coff[347 ] = 64'hffffef04ffff8122;
    assign coff[348 ] = 64'hffffeef8ffff8123;
    assign coff[349 ] = 64'hffffeeebffff8125;
    assign coff[350 ] = 64'hffffeedfffff8127;
    assign coff[351 ] = 64'hffffeed3ffff8128;
    assign coff[352 ] = 64'hffffeec6ffff812a;
    assign coff[353 ] = 64'hffffeebaffff812c;
    assign coff[354 ] = 64'hffffeeadffff812d;
    assign coff[355 ] = 64'hffffeea1ffff812f;
    assign coff[356 ] = 64'hffffee94ffff8131;
    assign coff[357 ] = 64'hffffee88ffff8133;
    assign coff[358 ] = 64'hffffee7bffff8134;
    assign coff[359 ] = 64'hffffee6fffff8136;
    assign coff[360 ] = 64'hffffee62ffff8138;
    assign coff[361 ] = 64'hffffee56ffff813a;
    assign coff[362 ] = 64'hffffee4affff813b;
    assign coff[363 ] = 64'hffffee3dffff813d;
    assign coff[364 ] = 64'hffffee31ffff813f;
    assign coff[365 ] = 64'hffffee24ffff8140;
    assign coff[366 ] = 64'hffffee18ffff8142;
    assign coff[367 ] = 64'hffffee0bffff8144;
    assign coff[368 ] = 64'hffffedffffff8146;
    assign coff[369 ] = 64'hffffedf2ffff8148;
    assign coff[370 ] = 64'hffffede6ffff8149;
    assign coff[371 ] = 64'hffffeddaffff814b;
    assign coff[372 ] = 64'hffffedcdffff814d;
    assign coff[373 ] = 64'hffffedc1ffff814f;
    assign coff[374 ] = 64'hffffedb4ffff8150;
    assign coff[375 ] = 64'hffffeda8ffff8152;
    assign coff[376 ] = 64'hffffed9bffff8154;
    assign coff[377 ] = 64'hffffed8fffff8156;
    assign coff[378 ] = 64'hffffed83ffff8158;
    assign coff[379 ] = 64'hffffed76ffff815a;
    assign coff[380 ] = 64'hffffed6affff815b;
    assign coff[381 ] = 64'hffffed5dffff815d;
    assign coff[382 ] = 64'hffffed51ffff815f;
    assign coff[383 ] = 64'hffffed44ffff8161;
    assign coff[384 ] = 64'hffffed38ffff8163;
    assign coff[385 ] = 64'hffffed2cffff8165;
    assign coff[386 ] = 64'hffffed1fffff8166;
    assign coff[387 ] = 64'hffffed13ffff8168;
    assign coff[388 ] = 64'hffffed06ffff816a;
    assign coff[389 ] = 64'hffffecfaffff816c;
    assign coff[390 ] = 64'hffffecedffff816e;
    assign coff[391 ] = 64'hffffece1ffff8170;
    assign coff[392 ] = 64'hffffecd5ffff8172;
    assign coff[393 ] = 64'hffffecc8ffff8173;
    assign coff[394 ] = 64'hffffecbcffff8175;
    assign coff[395 ] = 64'hffffecafffff8177;
    assign coff[396 ] = 64'hffffeca3ffff8179;
    assign coff[397 ] = 64'hffffec96ffff817b;
    assign coff[398 ] = 64'hffffec8affff817d;
    assign coff[399 ] = 64'hffffec7effff817f;
    assign coff[400 ] = 64'hffffec71ffff8181;
    assign coff[401 ] = 64'hffffec65ffff8183;
    assign coff[402 ] = 64'hffffec58ffff8185;
    assign coff[403 ] = 64'hffffec4cffff8187;
    assign coff[404 ] = 64'hffffec3fffff8188;
    assign coff[405 ] = 64'hffffec33ffff818a;
    assign coff[406 ] = 64'hffffec27ffff818c;
    assign coff[407 ] = 64'hffffec1affff818e;
    assign coff[408 ] = 64'hffffec0effff8190;
    assign coff[409 ] = 64'hffffec01ffff8192;
    assign coff[410 ] = 64'hffffebf5ffff8194;
    assign coff[411 ] = 64'hffffebe9ffff8196;
    assign coff[412 ] = 64'hffffebdcffff8198;
    assign coff[413 ] = 64'hffffebd0ffff819a;
    assign coff[414 ] = 64'hffffebc3ffff819c;
    assign coff[415 ] = 64'hffffebb7ffff819e;
    assign coff[416 ] = 64'hffffebabffff81a0;
    assign coff[417 ] = 64'hffffeb9effff81a2;
    assign coff[418 ] = 64'hffffeb92ffff81a4;
    assign coff[419 ] = 64'hffffeb85ffff81a6;
    assign coff[420 ] = 64'hffffeb79ffff81a8;
    assign coff[421 ] = 64'hffffeb6dffff81aa;
    assign coff[422 ] = 64'hffffeb60ffff81ac;
    assign coff[423 ] = 64'hffffeb54ffff81ae;
    assign coff[424 ] = 64'hffffeb47ffff81b0;
    assign coff[425 ] = 64'hffffeb3bffff81b2;
    assign coff[426 ] = 64'hffffeb2fffff81b4;
    assign coff[427 ] = 64'hffffeb22ffff81b6;
    assign coff[428 ] = 64'hffffeb16ffff81b8;
    assign coff[429 ] = 64'hffffeb09ffff81ba;
    assign coff[430 ] = 64'hffffeafdffff81bd;
    assign coff[431 ] = 64'hffffeaf1ffff81bf;
    assign coff[432 ] = 64'hffffeae4ffff81c1;
    assign coff[433 ] = 64'hffffead8ffff81c3;
    assign coff[434 ] = 64'hffffeacbffff81c5;
    assign coff[435 ] = 64'hffffeabfffff81c7;
    assign coff[436 ] = 64'hffffeab3ffff81c9;
    assign coff[437 ] = 64'hffffeaa6ffff81cb;
    assign coff[438 ] = 64'hffffea9affff81cd;
    assign coff[439 ] = 64'hffffea8dffff81cf;
    assign coff[440 ] = 64'hffffea81ffff81d1;
    assign coff[441 ] = 64'hffffea75ffff81d3;
    assign coff[442 ] = 64'hffffea68ffff81d6;
    assign coff[443 ] = 64'hffffea5cffff81d8;
    assign coff[444 ] = 64'hffffea4fffff81da;
    assign coff[445 ] = 64'hffffea43ffff81dc;
    assign coff[446 ] = 64'hffffea37ffff81de;
    assign coff[447 ] = 64'hffffea2affff81e0;
    assign coff[448 ] = 64'hffffea1effff81e2;
    assign coff[449 ] = 64'hffffea12ffff81e5;
    assign coff[450 ] = 64'hffffea05ffff81e7;
    assign coff[451 ] = 64'hffffe9f9ffff81e9;
    assign coff[452 ] = 64'hffffe9ecffff81eb;
    assign coff[453 ] = 64'hffffe9e0ffff81ed;
    assign coff[454 ] = 64'hffffe9d4ffff81ef;
    assign coff[455 ] = 64'hffffe9c7ffff81f2;
    assign coff[456 ] = 64'hffffe9bbffff81f4;
    assign coff[457 ] = 64'hffffe9afffff81f6;
    assign coff[458 ] = 64'hffffe9a2ffff81f8;
    assign coff[459 ] = 64'hffffe996ffff81fa;
    assign coff[460 ] = 64'hffffe989ffff81fd;
    assign coff[461 ] = 64'hffffe97dffff81ff;
    assign coff[462 ] = 64'hffffe971ffff8201;
    assign coff[463 ] = 64'hffffe964ffff8203;
    assign coff[464 ] = 64'hffffe958ffff8205;
    assign coff[465 ] = 64'hffffe94cffff8208;
    assign coff[466 ] = 64'hffffe93fffff820a;
    assign coff[467 ] = 64'hffffe933ffff820c;
    assign coff[468 ] = 64'hffffe926ffff820e;
    assign coff[469 ] = 64'hffffe91affff8211;
    assign coff[470 ] = 64'hffffe90effff8213;
    assign coff[471 ] = 64'hffffe901ffff8215;
    assign coff[472 ] = 64'hffffe8f5ffff8217;
    assign coff[473 ] = 64'hffffe8e9ffff821a;
    assign coff[474 ] = 64'hffffe8dcffff821c;
    assign coff[475 ] = 64'hffffe8d0ffff821e;
    assign coff[476 ] = 64'hffffe8c4ffff8220;
    assign coff[477 ] = 64'hffffe8b7ffff8223;
    assign coff[478 ] = 64'hffffe8abffff8225;
    assign coff[479 ] = 64'hffffe89fffff8227;
    assign coff[480 ] = 64'hffffe892ffff822a;
    assign coff[481 ] = 64'hffffe886ffff822c;
    assign coff[482 ] = 64'hffffe879ffff822e;
    assign coff[483 ] = 64'hffffe86dffff8231;
    assign coff[484 ] = 64'hffffe861ffff8233;
    assign coff[485 ] = 64'hffffe854ffff8235;
    assign coff[486 ] = 64'hffffe848ffff8237;
    assign coff[487 ] = 64'hffffe83cffff823a;
    assign coff[488 ] = 64'hffffe82fffff823c;
    assign coff[489 ] = 64'hffffe823ffff823e;
    assign coff[490 ] = 64'hffffe817ffff8241;
    assign coff[491 ] = 64'hffffe80affff8243;
    assign coff[492 ] = 64'hffffe7feffff8246;
    assign coff[493 ] = 64'hffffe7f2ffff8248;
    assign coff[494 ] = 64'hffffe7e5ffff824a;
    assign coff[495 ] = 64'hffffe7d9ffff824d;
    assign coff[496 ] = 64'hffffe7cdffff824f;
    assign coff[497 ] = 64'hffffe7c0ffff8251;
    assign coff[498 ] = 64'hffffe7b4ffff8254;
    assign coff[499 ] = 64'hffffe7a8ffff8256;
    assign coff[500 ] = 64'hffffe79bffff8259;
    assign coff[501 ] = 64'hffffe78fffff825b;
    assign coff[502 ] = 64'hffffe783ffff825d;
    assign coff[503 ] = 64'hffffe776ffff8260;
    assign coff[504 ] = 64'hffffe76affff8262;
    assign coff[505 ] = 64'hffffe75effff8265;
    assign coff[506 ] = 64'hffffe751ffff8267;
    assign coff[507 ] = 64'hffffe745ffff8269;
    assign coff[508 ] = 64'hffffe739ffff826c;
    assign coff[509 ] = 64'hffffe72cffff826e;
    assign coff[510 ] = 64'hffffe720ffff8271;
    assign coff[511 ] = 64'hffffe714ffff8273;
    assign coff[512 ] = 64'hffffe707ffff8276;
    assign coff[513 ] = 64'hffffe6fbffff8278;
    assign coff[514 ] = 64'hffffe6efffff827b;
    assign coff[515 ] = 64'hffffe6e2ffff827d;
    assign coff[516 ] = 64'hffffe6d6ffff827f;
    assign coff[517 ] = 64'hffffe6caffff8282;
    assign coff[518 ] = 64'hffffe6bdffff8284;
    assign coff[519 ] = 64'hffffe6b1ffff8287;
    assign coff[520 ] = 64'hffffe6a5ffff8289;
    assign coff[521 ] = 64'hffffe698ffff828c;
    assign coff[522 ] = 64'hffffe68cffff828e;
    assign coff[523 ] = 64'hffffe680ffff8291;
    assign coff[524 ] = 64'hffffe673ffff8293;
    assign coff[525 ] = 64'hffffe667ffff8296;
    assign coff[526 ] = 64'hffffe65bffff8298;
    assign coff[527 ] = 64'hffffe64fffff829b;
    assign coff[528 ] = 64'hffffe642ffff829d;
    assign coff[529 ] = 64'hffffe636ffff82a0;
    assign coff[530 ] = 64'hffffe62affff82a3;
    assign coff[531 ] = 64'hffffe61dffff82a5;
    assign coff[532 ] = 64'hffffe611ffff82a8;
    assign coff[533 ] = 64'hffffe605ffff82aa;
    assign coff[534 ] = 64'hffffe5f8ffff82ad;
    assign coff[535 ] = 64'hffffe5ecffff82af;
    assign coff[536 ] = 64'hffffe5e0ffff82b2;
    assign coff[537 ] = 64'hffffe5d3ffff82b4;
    assign coff[538 ] = 64'hffffe5c7ffff82b7;
    assign coff[539 ] = 64'hffffe5bbffff82ba;
    assign coff[540 ] = 64'hffffe5afffff82bc;
    assign coff[541 ] = 64'hffffe5a2ffff82bf;
    assign coff[542 ] = 64'hffffe596ffff82c1;
    assign coff[543 ] = 64'hffffe58affff82c4;
    assign coff[544 ] = 64'hffffe57dffff82c6;
    assign coff[545 ] = 64'hffffe571ffff82c9;
    assign coff[546 ] = 64'hffffe565ffff82cc;
    assign coff[547 ] = 64'hffffe558ffff82ce;
    assign coff[548 ] = 64'hffffe54cffff82d1;
    assign coff[549 ] = 64'hffffe540ffff82d4;
    assign coff[550 ] = 64'hffffe534ffff82d6;
    assign coff[551 ] = 64'hffffe527ffff82d9;
    assign coff[552 ] = 64'hffffe51bffff82db;
    assign coff[553 ] = 64'hffffe50fffff82de;
    assign coff[554 ] = 64'hffffe502ffff82e1;
    assign coff[555 ] = 64'hffffe4f6ffff82e3;
    assign coff[556 ] = 64'hffffe4eaffff82e6;
    assign coff[557 ] = 64'hffffe4deffff82e9;
    assign coff[558 ] = 64'hffffe4d1ffff82eb;
    assign coff[559 ] = 64'hffffe4c5ffff82ee;
    assign coff[560 ] = 64'hffffe4b9ffff82f1;
    assign coff[561 ] = 64'hffffe4adffff82f3;
    assign coff[562 ] = 64'hffffe4a0ffff82f6;
    assign coff[563 ] = 64'hffffe494ffff82f9;
    assign coff[564 ] = 64'hffffe488ffff82fb;
    assign coff[565 ] = 64'hffffe47bffff82fe;
    assign coff[566 ] = 64'hffffe46fffff8301;
    assign coff[567 ] = 64'hffffe463ffff8304;
    assign coff[568 ] = 64'hffffe457ffff8306;
    assign coff[569 ] = 64'hffffe44affff8309;
    assign coff[570 ] = 64'hffffe43effff830c;
    assign coff[571 ] = 64'hffffe432ffff830e;
    assign coff[572 ] = 64'hffffe426ffff8311;
    assign coff[573 ] = 64'hffffe419ffff8314;
    assign coff[574 ] = 64'hffffe40dffff8317;
    assign coff[575 ] = 64'hffffe401ffff8319;
    assign coff[576 ] = 64'hffffe3f4ffff831c;
    assign coff[577 ] = 64'hffffe3e8ffff831f;
    assign coff[578 ] = 64'hffffe3dcffff8322;
    assign coff[579 ] = 64'hffffe3d0ffff8324;
    assign coff[580 ] = 64'hffffe3c3ffff8327;
    assign coff[581 ] = 64'hffffe3b7ffff832a;
    assign coff[582 ] = 64'hffffe3abffff832d;
    assign coff[583 ] = 64'hffffe39fffff8330;
    assign coff[584 ] = 64'hffffe392ffff8332;
    assign coff[585 ] = 64'hffffe386ffff8335;
    assign coff[586 ] = 64'hffffe37affff8338;
    assign coff[587 ] = 64'hffffe36effff833b;
    assign coff[588 ] = 64'hffffe361ffff833e;
    assign coff[589 ] = 64'hffffe355ffff8340;
    assign coff[590 ] = 64'hffffe349ffff8343;
    assign coff[591 ] = 64'hffffe33dffff8346;
    assign coff[592 ] = 64'hffffe330ffff8349;
    assign coff[593 ] = 64'hffffe324ffff834c;
    assign coff[594 ] = 64'hffffe318ffff834f;
    assign coff[595 ] = 64'hffffe30cffff8351;
    assign coff[596 ] = 64'hffffe2ffffff8354;
    assign coff[597 ] = 64'hffffe2f3ffff8357;
    assign coff[598 ] = 64'hffffe2e7ffff835a;
    assign coff[599 ] = 64'hffffe2dbffff835d;
    assign coff[600 ] = 64'hffffe2cfffff8360;
    assign coff[601 ] = 64'hffffe2c2ffff8362;
    assign coff[602 ] = 64'hffffe2b6ffff8365;
    assign coff[603 ] = 64'hffffe2aaffff8368;
    assign coff[604 ] = 64'hffffe29effff836b;
    assign coff[605 ] = 64'hffffe291ffff836e;
    assign coff[606 ] = 64'hffffe285ffff8371;
    assign coff[607 ] = 64'hffffe279ffff8374;
    assign coff[608 ] = 64'hffffe26dffff8377;
    assign coff[609 ] = 64'hffffe260ffff837a;
    assign coff[610 ] = 64'hffffe254ffff837d;
    assign coff[611 ] = 64'hffffe248ffff837f;
    assign coff[612 ] = 64'hffffe23cffff8382;
    assign coff[613 ] = 64'hffffe230ffff8385;
    assign coff[614 ] = 64'hffffe223ffff8388;
    assign coff[615 ] = 64'hffffe217ffff838b;
    assign coff[616 ] = 64'hffffe20bffff838e;
    assign coff[617 ] = 64'hffffe1ffffff8391;
    assign coff[618 ] = 64'hffffe1f2ffff8394;
    assign coff[619 ] = 64'hffffe1e6ffff8397;
    assign coff[620 ] = 64'hffffe1daffff839a;
    assign coff[621 ] = 64'hffffe1ceffff839d;
    assign coff[622 ] = 64'hffffe1c2ffff83a0;
    assign coff[623 ] = 64'hffffe1b5ffff83a3;
    assign coff[624 ] = 64'hffffe1a9ffff83a6;
    assign coff[625 ] = 64'hffffe19dffff83a9;
    assign coff[626 ] = 64'hffffe191ffff83ac;
    assign coff[627 ] = 64'hffffe185ffff83af;
    assign coff[628 ] = 64'hffffe178ffff83b2;
    assign coff[629 ] = 64'hffffe16cffff83b5;
    assign coff[630 ] = 64'hffffe160ffff83b8;
    assign coff[631 ] = 64'hffffe154ffff83bb;
    assign coff[632 ] = 64'hffffe148ffff83be;
    assign coff[633 ] = 64'hffffe13bffff83c1;
    assign coff[634 ] = 64'hffffe12fffff83c4;
    assign coff[635 ] = 64'hffffe123ffff83c7;
    assign coff[636 ] = 64'hffffe117ffff83ca;
    assign coff[637 ] = 64'hffffe10bffff83cd;
    assign coff[638 ] = 64'hffffe0feffff83d0;
    assign coff[639 ] = 64'hffffe0f2ffff83d3;
    assign coff[640 ] = 64'hffffe0e6ffff83d6;
    assign coff[641 ] = 64'hffffe0daffff83d9;
    assign coff[642 ] = 64'hffffe0ceffff83dc;
    assign coff[643 ] = 64'hffffe0c1ffff83df;
    assign coff[644 ] = 64'hffffe0b5ffff83e2;
    assign coff[645 ] = 64'hffffe0a9ffff83e5;
    assign coff[646 ] = 64'hffffe09dffff83e8;
    assign coff[647 ] = 64'hffffe091ffff83ec;
    assign coff[648 ] = 64'hffffe085ffff83ef;
    assign coff[649 ] = 64'hffffe078ffff83f2;
    assign coff[650 ] = 64'hffffe06cffff83f5;
    assign coff[651 ] = 64'hffffe060ffff83f8;
    assign coff[652 ] = 64'hffffe054ffff83fb;
    assign coff[653 ] = 64'hffffe048ffff83fe;
    assign coff[654 ] = 64'hffffe03bffff8401;
    assign coff[655 ] = 64'hffffe02fffff8404;
    assign coff[656 ] = 64'hffffe023ffff8407;
    assign coff[657 ] = 64'hffffe017ffff840b;
    assign coff[658 ] = 64'hffffe00bffff840e;
    assign coff[659 ] = 64'hffffdfffffff8411;
    assign coff[660 ] = 64'hffffdff2ffff8414;
    assign coff[661 ] = 64'hffffdfe6ffff8417;
    assign coff[662 ] = 64'hffffdfdaffff841a;
    assign coff[663 ] = 64'hffffdfceffff841d;
    assign coff[664 ] = 64'hffffdfc2ffff8421;
    assign coff[665 ] = 64'hffffdfb6ffff8424;
    assign coff[666 ] = 64'hffffdfa9ffff8427;
    assign coff[667 ] = 64'hffffdf9dffff842a;
    assign coff[668 ] = 64'hffffdf91ffff842d;
    assign coff[669 ] = 64'hffffdf85ffff8431;
    assign coff[670 ] = 64'hffffdf79ffff8434;
    assign coff[671 ] = 64'hffffdf6dffff8437;
    assign coff[672 ] = 64'hffffdf61ffff843a;
    assign coff[673 ] = 64'hffffdf54ffff843d;
    assign coff[674 ] = 64'hffffdf48ffff8441;
    assign coff[675 ] = 64'hffffdf3cffff8444;
    assign coff[676 ] = 64'hffffdf30ffff8447;
    assign coff[677 ] = 64'hffffdf24ffff844a;
    assign coff[678 ] = 64'hffffdf18ffff844d;
    assign coff[679 ] = 64'hffffdf0cffff8451;
    assign coff[680 ] = 64'hffffdeffffff8454;
    assign coff[681 ] = 64'hffffdef3ffff8457;
    assign coff[682 ] = 64'hffffdee7ffff845a;
    assign coff[683 ] = 64'hffffdedbffff845e;
    assign coff[684 ] = 64'hffffdecfffff8461;
    assign coff[685 ] = 64'hffffdec3ffff8464;
    assign coff[686 ] = 64'hffffdeb7ffff8467;
    assign coff[687 ] = 64'hffffdeaaffff846b;
    assign coff[688 ] = 64'hffffde9effff846e;
    assign coff[689 ] = 64'hffffde92ffff8471;
    assign coff[690 ] = 64'hffffde86ffff8475;
    assign coff[691 ] = 64'hffffde7affff8478;
    assign coff[692 ] = 64'hffffde6effff847b;
    assign coff[693 ] = 64'hffffde62ffff847e;
    assign coff[694 ] = 64'hffffde56ffff8482;
    assign coff[695 ] = 64'hffffde49ffff8485;
    assign coff[696 ] = 64'hffffde3dffff8488;
    assign coff[697 ] = 64'hffffde31ffff848c;
    assign coff[698 ] = 64'hffffde25ffff848f;
    assign coff[699 ] = 64'hffffde19ffff8492;
    assign coff[700 ] = 64'hffffde0dffff8496;
    assign coff[701 ] = 64'hffffde01ffff8499;
    assign coff[702 ] = 64'hffffddf5ffff849c;
    assign coff[703 ] = 64'hffffdde8ffff84a0;
    assign coff[704 ] = 64'hffffdddcffff84a3;
    assign coff[705 ] = 64'hffffddd0ffff84a6;
    assign coff[706 ] = 64'hffffddc4ffff84aa;
    assign coff[707 ] = 64'hffffddb8ffff84ad;
    assign coff[708 ] = 64'hffffddacffff84b0;
    assign coff[709 ] = 64'hffffdda0ffff84b4;
    assign coff[710 ] = 64'hffffdd94ffff84b7;
    assign coff[711 ] = 64'hffffdd88ffff84bb;
    assign coff[712 ] = 64'hffffdd7cffff84be;
    assign coff[713 ] = 64'hffffdd6fffff84c1;
    assign coff[714 ] = 64'hffffdd63ffff84c5;
    assign coff[715 ] = 64'hffffdd57ffff84c8;
    assign coff[716 ] = 64'hffffdd4bffff84cc;
    assign coff[717 ] = 64'hffffdd3fffff84cf;
    assign coff[718 ] = 64'hffffdd33ffff84d2;
    assign coff[719 ] = 64'hffffdd27ffff84d6;
    assign coff[720 ] = 64'hffffdd1bffff84d9;
    assign coff[721 ] = 64'hffffdd0fffff84dd;
    assign coff[722 ] = 64'hffffdd03ffff84e0;
    assign coff[723 ] = 64'hffffdcf6ffff84e4;
    assign coff[724 ] = 64'hffffdceaffff84e7;
    assign coff[725 ] = 64'hffffdcdeffff84ea;
    assign coff[726 ] = 64'hffffdcd2ffff84ee;
    assign coff[727 ] = 64'hffffdcc6ffff84f1;
    assign coff[728 ] = 64'hffffdcbaffff84f5;
    assign coff[729 ] = 64'hffffdcaeffff84f8;
    assign coff[730 ] = 64'hffffdca2ffff84fc;
    assign coff[731 ] = 64'hffffdc96ffff84ff;
    assign coff[732 ] = 64'hffffdc8affff8503;
    assign coff[733 ] = 64'hffffdc7effff8506;
    assign coff[734 ] = 64'hffffdc72ffff850a;
    assign coff[735 ] = 64'hffffdc66ffff850d;
    assign coff[736 ] = 64'hffffdc59ffff8511;
    assign coff[737 ] = 64'hffffdc4dffff8514;
    assign coff[738 ] = 64'hffffdc41ffff8518;
    assign coff[739 ] = 64'hffffdc35ffff851b;
    assign coff[740 ] = 64'hffffdc29ffff851f;
    assign coff[741 ] = 64'hffffdc1dffff8522;
    assign coff[742 ] = 64'hffffdc11ffff8526;
    assign coff[743 ] = 64'hffffdc05ffff8529;
    assign coff[744 ] = 64'hffffdbf9ffff852d;
    assign coff[745 ] = 64'hffffdbedffff8530;
    assign coff[746 ] = 64'hffffdbe1ffff8534;
    assign coff[747 ] = 64'hffffdbd5ffff8537;
    assign coff[748 ] = 64'hffffdbc9ffff853b;
    assign coff[749 ] = 64'hffffdbbdffff853f;
    assign coff[750 ] = 64'hffffdbb1ffff8542;
    assign coff[751 ] = 64'hffffdba5ffff8546;
    assign coff[752 ] = 64'hffffdb99ffff8549;
    assign coff[753 ] = 64'hffffdb8cffff854d;
    assign coff[754 ] = 64'hffffdb80ffff8550;
    assign coff[755 ] = 64'hffffdb74ffff8554;
    assign coff[756 ] = 64'hffffdb68ffff8558;
    assign coff[757 ] = 64'hffffdb5cffff855b;
    assign coff[758 ] = 64'hffffdb50ffff855f;
    assign coff[759 ] = 64'hffffdb44ffff8562;
    assign coff[760 ] = 64'hffffdb38ffff8566;
    assign coff[761 ] = 64'hffffdb2cffff856a;
    assign coff[762 ] = 64'hffffdb20ffff856d;
    assign coff[763 ] = 64'hffffdb14ffff8571;
    assign coff[764 ] = 64'hffffdb08ffff8574;
    assign coff[765 ] = 64'hffffdafcffff8578;
    assign coff[766 ] = 64'hffffdaf0ffff857c;
    assign coff[767 ] = 64'hffffdae4ffff857f;
    assign coff[768 ] = 64'hffffdad8ffff8583;
    assign coff[769 ] = 64'hffffdaccffff8587;
    assign coff[770 ] = 64'hffffdac0ffff858a;
    assign coff[771 ] = 64'hffffdab4ffff858e;
    assign coff[772 ] = 64'hffffdaa8ffff8592;
    assign coff[773 ] = 64'hffffda9cffff8595;
    assign coff[774 ] = 64'hffffda90ffff8599;
    assign coff[775 ] = 64'hffffda84ffff859d;
    assign coff[776 ] = 64'hffffda78ffff85a0;
    assign coff[777 ] = 64'hffffda6cffff85a4;
    assign coff[778 ] = 64'hffffda60ffff85a8;
    assign coff[779 ] = 64'hffffda54ffff85ab;
    assign coff[780 ] = 64'hffffda48ffff85af;
    assign coff[781 ] = 64'hffffda3cffff85b3;
    assign coff[782 ] = 64'hffffda30ffff85b7;
    assign coff[783 ] = 64'hffffda24ffff85ba;
    assign coff[784 ] = 64'hffffda18ffff85be;
    assign coff[785 ] = 64'hffffda0cffff85c2;
    assign coff[786 ] = 64'hffffda00ffff85c5;
    assign coff[787 ] = 64'hffffd9f4ffff85c9;
    assign coff[788 ] = 64'hffffd9e8ffff85cd;
    assign coff[789 ] = 64'hffffd9dcffff85d1;
    assign coff[790 ] = 64'hffffd9d0ffff85d4;
    assign coff[791 ] = 64'hffffd9c4ffff85d8;
    assign coff[792 ] = 64'hffffd9b8ffff85dc;
    assign coff[793 ] = 64'hffffd9acffff85e0;
    assign coff[794 ] = 64'hffffd9a0ffff85e3;
    assign coff[795 ] = 64'hffffd994ffff85e7;
    assign coff[796 ] = 64'hffffd988ffff85eb;
    assign coff[797 ] = 64'hffffd97cffff85ef;
    assign coff[798 ] = 64'hffffd970ffff85f2;
    assign coff[799 ] = 64'hffffd964ffff85f6;
    assign coff[800 ] = 64'hffffd958ffff85fa;
    assign coff[801 ] = 64'hffffd94cffff85fe;
    assign coff[802 ] = 64'hffffd940ffff8602;
    assign coff[803 ] = 64'hffffd934ffff8605;
    assign coff[804 ] = 64'hffffd928ffff8609;
    assign coff[805 ] = 64'hffffd91cffff860d;
    assign coff[806 ] = 64'hffffd910ffff8611;
    assign coff[807 ] = 64'hffffd904ffff8615;
    assign coff[808 ] = 64'hffffd8f8ffff8619;
    assign coff[809 ] = 64'hffffd8ecffff861c;
    assign coff[810 ] = 64'hffffd8e0ffff8620;
    assign coff[811 ] = 64'hffffd8d4ffff8624;
    assign coff[812 ] = 64'hffffd8c8ffff8628;
    assign coff[813 ] = 64'hffffd8bcffff862c;
    assign coff[814 ] = 64'hffffd8b0ffff8630;
    assign coff[815 ] = 64'hffffd8a4ffff8634;
    assign coff[816 ] = 64'hffffd898ffff8637;
    assign coff[817 ] = 64'hffffd88cffff863b;
    assign coff[818 ] = 64'hffffd880ffff863f;
    assign coff[819 ] = 64'hffffd875ffff8643;
    assign coff[820 ] = 64'hffffd869ffff8647;
    assign coff[821 ] = 64'hffffd85dffff864b;
    assign coff[822 ] = 64'hffffd851ffff864f;
    assign coff[823 ] = 64'hffffd845ffff8653;
    assign coff[824 ] = 64'hffffd839ffff8656;
    assign coff[825 ] = 64'hffffd82dffff865a;
    assign coff[826 ] = 64'hffffd821ffff865e;
    assign coff[827 ] = 64'hffffd815ffff8662;
    assign coff[828 ] = 64'hffffd809ffff8666;
    assign coff[829 ] = 64'hffffd7fdffff866a;
    assign coff[830 ] = 64'hffffd7f1ffff866e;
    assign coff[831 ] = 64'hffffd7e5ffff8672;
    assign coff[832 ] = 64'hffffd7d9ffff8676;
    assign coff[833 ] = 64'hffffd7cdffff867a;
    assign coff[834 ] = 64'hffffd7c1ffff867e;
    assign coff[835 ] = 64'hffffd7b5ffff8682;
    assign coff[836 ] = 64'hffffd7aaffff8686;
    assign coff[837 ] = 64'hffffd79effff868a;
    assign coff[838 ] = 64'hffffd792ffff868e;
    assign coff[839 ] = 64'hffffd786ffff8692;
    assign coff[840 ] = 64'hffffd77affff8696;
    assign coff[841 ] = 64'hffffd76effff869a;
    assign coff[842 ] = 64'hffffd762ffff869e;
    assign coff[843 ] = 64'hffffd756ffff86a1;
    assign coff[844 ] = 64'hffffd74affff86a5;
    assign coff[845 ] = 64'hffffd73effff86a9;
    assign coff[846 ] = 64'hffffd732ffff86ad;
    assign coff[847 ] = 64'hffffd726ffff86b2;
    assign coff[848 ] = 64'hffffd71bffff86b6;
    assign coff[849 ] = 64'hffffd70fffff86ba;
    assign coff[850 ] = 64'hffffd703ffff86be;
    assign coff[851 ] = 64'hffffd6f7ffff86c2;
    assign coff[852 ] = 64'hffffd6ebffff86c6;
    assign coff[853 ] = 64'hffffd6dfffff86ca;
    assign coff[854 ] = 64'hffffd6d3ffff86ce;
    assign coff[855 ] = 64'hffffd6c7ffff86d2;
    assign coff[856 ] = 64'hffffd6bbffff86d6;
    assign coff[857 ] = 64'hffffd6afffff86da;
    assign coff[858 ] = 64'hffffd6a4ffff86de;
    assign coff[859 ] = 64'hffffd698ffff86e2;
    assign coff[860 ] = 64'hffffd68cffff86e6;
    assign coff[861 ] = 64'hffffd680ffff86ea;
    assign coff[862 ] = 64'hffffd674ffff86ee;
    assign coff[863 ] = 64'hffffd668ffff86f2;
    assign coff[864 ] = 64'hffffd65cffff86f6;
    assign coff[865 ] = 64'hffffd650ffff86fa;
    assign coff[866 ] = 64'hffffd644ffff86ff;
    assign coff[867 ] = 64'hffffd639ffff8703;
    assign coff[868 ] = 64'hffffd62dffff8707;
    assign coff[869 ] = 64'hffffd621ffff870b;
    assign coff[870 ] = 64'hffffd615ffff870f;
    assign coff[871 ] = 64'hffffd609ffff8713;
    assign coff[872 ] = 64'hffffd5fdffff8717;
    assign coff[873 ] = 64'hffffd5f1ffff871b;
    assign coff[874 ] = 64'hffffd5e5ffff871f;
    assign coff[875 ] = 64'hffffd5daffff8724;
    assign coff[876 ] = 64'hffffd5ceffff8728;
    assign coff[877 ] = 64'hffffd5c2ffff872c;
    assign coff[878 ] = 64'hffffd5b6ffff8730;
    assign coff[879 ] = 64'hffffd5aaffff8734;
    assign coff[880 ] = 64'hffffd59effff8738;
    assign coff[881 ] = 64'hffffd592ffff873c;
    assign coff[882 ] = 64'hffffd587ffff8741;
    assign coff[883 ] = 64'hffffd57bffff8745;
    assign coff[884 ] = 64'hffffd56fffff8749;
    assign coff[885 ] = 64'hffffd563ffff874d;
    assign coff[886 ] = 64'hffffd557ffff8751;
    assign coff[887 ] = 64'hffffd54bffff8756;
    assign coff[888 ] = 64'hffffd53fffff875a;
    assign coff[889 ] = 64'hffffd534ffff875e;
    assign coff[890 ] = 64'hffffd528ffff8762;
    assign coff[891 ] = 64'hffffd51cffff8766;
    assign coff[892 ] = 64'hffffd510ffff876b;
    assign coff[893 ] = 64'hffffd504ffff876f;
    assign coff[894 ] = 64'hffffd4f8ffff8773;
    assign coff[895 ] = 64'hffffd4edffff8777;
    assign coff[896 ] = 64'hffffd4e1ffff877b;
    assign coff[897 ] = 64'hffffd4d5ffff8780;
    assign coff[898 ] = 64'hffffd4c9ffff8784;
    assign coff[899 ] = 64'hffffd4bdffff8788;
    assign coff[900 ] = 64'hffffd4b1ffff878c;
    assign coff[901 ] = 64'hffffd4a6ffff8791;
    assign coff[902 ] = 64'hffffd49affff8795;
    assign coff[903 ] = 64'hffffd48effff8799;
    assign coff[904 ] = 64'hffffd482ffff879d;
    assign coff[905 ] = 64'hffffd476ffff87a2;
    assign coff[906 ] = 64'hffffd46bffff87a6;
    assign coff[907 ] = 64'hffffd45fffff87aa;
    assign coff[908 ] = 64'hffffd453ffff87af;
    assign coff[909 ] = 64'hffffd447ffff87b3;
    assign coff[910 ] = 64'hffffd43bffff87b7;
    assign coff[911 ] = 64'hffffd430ffff87bb;
    assign coff[912 ] = 64'hffffd424ffff87c0;
    assign coff[913 ] = 64'hffffd418ffff87c4;
    assign coff[914 ] = 64'hffffd40cffff87c8;
    assign coff[915 ] = 64'hffffd400ffff87cd;
    assign coff[916 ] = 64'hffffd3f4ffff87d1;
    assign coff[917 ] = 64'hffffd3e9ffff87d5;
    assign coff[918 ] = 64'hffffd3ddffff87da;
    assign coff[919 ] = 64'hffffd3d1ffff87de;
    assign coff[920 ] = 64'hffffd3c5ffff87e2;
    assign coff[921 ] = 64'hffffd3baffff87e7;
    assign coff[922 ] = 64'hffffd3aeffff87eb;
    assign coff[923 ] = 64'hffffd3a2ffff87ef;
    assign coff[924 ] = 64'hffffd396ffff87f4;
    assign coff[925 ] = 64'hffffd38affff87f8;
    assign coff[926 ] = 64'hffffd37fffff87fd;
    assign coff[927 ] = 64'hffffd373ffff8801;
    assign coff[928 ] = 64'hffffd367ffff8805;
    assign coff[929 ] = 64'hffffd35bffff880a;
    assign coff[930 ] = 64'hffffd34fffff880e;
    assign coff[931 ] = 64'hffffd344ffff8812;
    assign coff[932 ] = 64'hffffd338ffff8817;
    assign coff[933 ] = 64'hffffd32cffff881b;
    assign coff[934 ] = 64'hffffd320ffff8820;
    assign coff[935 ] = 64'hffffd315ffff8824;
    assign coff[936 ] = 64'hffffd309ffff8828;
    assign coff[937 ] = 64'hffffd2fdffff882d;
    assign coff[938 ] = 64'hffffd2f1ffff8831;
    assign coff[939 ] = 64'hffffd2e6ffff8836;
    assign coff[940 ] = 64'hffffd2daffff883a;
    assign coff[941 ] = 64'hffffd2ceffff883f;
    assign coff[942 ] = 64'hffffd2c2ffff8843;
    assign coff[943 ] = 64'hffffd2b7ffff8847;
    assign coff[944 ] = 64'hffffd2abffff884c;
    assign coff[945 ] = 64'hffffd29fffff8850;
    assign coff[946 ] = 64'hffffd293ffff8855;
    assign coff[947 ] = 64'hffffd288ffff8859;
    assign coff[948 ] = 64'hffffd27cffff885e;
    assign coff[949 ] = 64'hffffd270ffff8862;
    assign coff[950 ] = 64'hffffd264ffff8867;
    assign coff[951 ] = 64'hffffd259ffff886b;
    assign coff[952 ] = 64'hffffd24dffff8870;
    assign coff[953 ] = 64'hffffd241ffff8874;
    assign coff[954 ] = 64'hffffd235ffff8879;
    assign coff[955 ] = 64'hffffd22affff887d;
    assign coff[956 ] = 64'hffffd21effff8882;
    assign coff[957 ] = 64'hffffd212ffff8886;
    assign coff[958 ] = 64'hffffd206ffff888b;
    assign coff[959 ] = 64'hffffd1fbffff888f;
    assign coff[960 ] = 64'hffffd1efffff8894;
    assign coff[961 ] = 64'hffffd1e3ffff8898;
    assign coff[962 ] = 64'hffffd1d8ffff889d;
    assign coff[963 ] = 64'hffffd1ccffff88a1;
    assign coff[964 ] = 64'hffffd1c0ffff88a6;
    assign coff[965 ] = 64'hffffd1b4ffff88aa;
    assign coff[966 ] = 64'hffffd1a9ffff88af;
    assign coff[967 ] = 64'hffffd19dffff88b3;
    assign coff[968 ] = 64'hffffd191ffff88b8;
    assign coff[969 ] = 64'hffffd186ffff88bd;
    assign coff[970 ] = 64'hffffd17affff88c1;
    assign coff[971 ] = 64'hffffd16effff88c6;
    assign coff[972 ] = 64'hffffd162ffff88ca;
    assign coff[973 ] = 64'hffffd157ffff88cf;
    assign coff[974 ] = 64'hffffd14bffff88d3;
    assign coff[975 ] = 64'hffffd13fffff88d8;
    assign coff[976 ] = 64'hffffd134ffff88dd;
    assign coff[977 ] = 64'hffffd128ffff88e1;
    assign coff[978 ] = 64'hffffd11cffff88e6;
    assign coff[979 ] = 64'hffffd111ffff88ea;
    assign coff[980 ] = 64'hffffd105ffff88ef;
    assign coff[981 ] = 64'hffffd0f9ffff88f4;
    assign coff[982 ] = 64'hffffd0edffff88f8;
    assign coff[983 ] = 64'hffffd0e2ffff88fd;
    assign coff[984 ] = 64'hffffd0d6ffff8902;
    assign coff[985 ] = 64'hffffd0caffff8906;
    assign coff[986 ] = 64'hffffd0bfffff890b;
    assign coff[987 ] = 64'hffffd0b3ffff890f;
    assign coff[988 ] = 64'hffffd0a7ffff8914;
    assign coff[989 ] = 64'hffffd09cffff8919;
    assign coff[990 ] = 64'hffffd090ffff891d;
    assign coff[991 ] = 64'hffffd084ffff8922;
    assign coff[992 ] = 64'hffffd079ffff8927;
    assign coff[993 ] = 64'hffffd06dffff892b;
    assign coff[994 ] = 64'hffffd061ffff8930;
    assign coff[995 ] = 64'hffffd056ffff8935;
    assign coff[996 ] = 64'hffffd04affff8939;
    assign coff[997 ] = 64'hffffd03effff893e;
    assign coff[998 ] = 64'hffffd033ffff8943;
    assign coff[999 ] = 64'hffffd027ffff8947;
    assign coff[1000] = 64'hffffd01bffff894c;
    assign coff[1001] = 64'hffffd010ffff8951;
    assign coff[1002] = 64'hffffd004ffff8956;
    assign coff[1003] = 64'hffffcff8ffff895a;
    assign coff[1004] = 64'hffffcfedffff895f;
    assign coff[1005] = 64'hffffcfe1ffff8964;
    assign coff[1006] = 64'hffffcfd6ffff8968;
    assign coff[1007] = 64'hffffcfcaffff896d;
    assign coff[1008] = 64'hffffcfbeffff8972;
    assign coff[1009] = 64'hffffcfb3ffff8977;
    assign coff[1010] = 64'hffffcfa7ffff897b;
    assign coff[1011] = 64'hffffcf9bffff8980;
    assign coff[1012] = 64'hffffcf90ffff8985;
    assign coff[1013] = 64'hffffcf84ffff898a;
    assign coff[1014] = 64'hffffcf78ffff898e;
    assign coff[1015] = 64'hffffcf6dffff8993;
    assign coff[1016] = 64'hffffcf61ffff8998;
    assign coff[1017] = 64'hffffcf56ffff899d;
    assign coff[1018] = 64'hffffcf4affff89a2;
    assign coff[1019] = 64'hffffcf3effff89a6;
    assign coff[1020] = 64'hffffcf33ffff89ab;
    assign coff[1021] = 64'hffffcf27ffff89b0;
    assign coff[1022] = 64'hffffcf1bffff89b5;
    assign coff[1023] = 64'hffffcf10ffff89ba;
    assign coff[1024] = 64'hffffcf04ffff89be;
    assign coff[1025] = 64'hffffcef9ffff89c3;
    assign coff[1026] = 64'hffffceedffff89c8;
    assign coff[1027] = 64'hffffcee1ffff89cd;
    assign coff[1028] = 64'hffffced6ffff89d2;
    assign coff[1029] = 64'hffffcecaffff89d6;
    assign coff[1030] = 64'hffffcebfffff89db;
    assign coff[1031] = 64'hffffceb3ffff89e0;
    assign coff[1032] = 64'hffffcea7ffff89e5;
    assign coff[1033] = 64'hffffce9cffff89ea;
    assign coff[1034] = 64'hffffce90ffff89ef;
    assign coff[1035] = 64'hffffce85ffff89f3;
    assign coff[1036] = 64'hffffce79ffff89f8;
    assign coff[1037] = 64'hffffce6dffff89fd;
    assign coff[1038] = 64'hffffce62ffff8a02;
    assign coff[1039] = 64'hffffce56ffff8a07;
    assign coff[1040] = 64'hffffce4bffff8a0c;
    assign coff[1041] = 64'hffffce3fffff8a11;
    assign coff[1042] = 64'hffffce34ffff8a16;
    assign coff[1043] = 64'hffffce28ffff8a1a;
    assign coff[1044] = 64'hffffce1cffff8a1f;
    assign coff[1045] = 64'hffffce11ffff8a24;
    assign coff[1046] = 64'hffffce05ffff8a29;
    assign coff[1047] = 64'hffffcdfaffff8a2e;
    assign coff[1048] = 64'hffffcdeeffff8a33;
    assign coff[1049] = 64'hffffcde3ffff8a38;
    assign coff[1050] = 64'hffffcdd7ffff8a3d;
    assign coff[1051] = 64'hffffcdcbffff8a42;
    assign coff[1052] = 64'hffffcdc0ffff8a47;
    assign coff[1053] = 64'hffffcdb4ffff8a4c;
    assign coff[1054] = 64'hffffcda9ffff8a51;
    assign coff[1055] = 64'hffffcd9dffff8a56;
    assign coff[1056] = 64'hffffcd92ffff8a5a;
    assign coff[1057] = 64'hffffcd86ffff8a5f;
    assign coff[1058] = 64'hffffcd7bffff8a64;
    assign coff[1059] = 64'hffffcd6fffff8a69;
    assign coff[1060] = 64'hffffcd63ffff8a6e;
    assign coff[1061] = 64'hffffcd58ffff8a73;
    assign coff[1062] = 64'hffffcd4cffff8a78;
    assign coff[1063] = 64'hffffcd41ffff8a7d;
    assign coff[1064] = 64'hffffcd35ffff8a82;
    assign coff[1065] = 64'hffffcd2affff8a87;
    assign coff[1066] = 64'hffffcd1effff8a8c;
    assign coff[1067] = 64'hffffcd13ffff8a91;
    assign coff[1068] = 64'hffffcd07ffff8a96;
    assign coff[1069] = 64'hffffccfcffff8a9b;
    assign coff[1070] = 64'hffffccf0ffff8aa0;
    assign coff[1071] = 64'hffffcce5ffff8aa5;
    assign coff[1072] = 64'hffffccd9ffff8aaa;
    assign coff[1073] = 64'hffffccceffff8aaf;
    assign coff[1074] = 64'hffffccc2ffff8ab4;
    assign coff[1075] = 64'hffffccb7ffff8ab9;
    assign coff[1076] = 64'hffffccabffff8abe;
    assign coff[1077] = 64'hffffcca0ffff8ac3;
    assign coff[1078] = 64'hffffcc94ffff8ac8;
    assign coff[1079] = 64'hffffcc89ffff8ace;
    assign coff[1080] = 64'hffffcc7dffff8ad3;
    assign coff[1081] = 64'hffffcc72ffff8ad8;
    assign coff[1082] = 64'hffffcc66ffff8add;
    assign coff[1083] = 64'hffffcc5bffff8ae2;
    assign coff[1084] = 64'hffffcc4fffff8ae7;
    assign coff[1085] = 64'hffffcc44ffff8aec;
    assign coff[1086] = 64'hffffcc38ffff8af1;
    assign coff[1087] = 64'hffffcc2dffff8af6;
    assign coff[1088] = 64'hffffcc21ffff8afb;
    assign coff[1089] = 64'hffffcc16ffff8b00;
    assign coff[1090] = 64'hffffcc0affff8b05;
    assign coff[1091] = 64'hffffcbffffff8b0a;
    assign coff[1092] = 64'hffffcbf3ffff8b10;
    assign coff[1093] = 64'hffffcbe8ffff8b15;
    assign coff[1094] = 64'hffffcbdcffff8b1a;
    assign coff[1095] = 64'hffffcbd1ffff8b1f;
    assign coff[1096] = 64'hffffcbc5ffff8b24;
    assign coff[1097] = 64'hffffcbbaffff8b29;
    assign coff[1098] = 64'hffffcbaeffff8b2e;
    assign coff[1099] = 64'hffffcba3ffff8b33;
    assign coff[1100] = 64'hffffcb97ffff8b39;
    assign coff[1101] = 64'hffffcb8cffff8b3e;
    assign coff[1102] = 64'hffffcb80ffff8b43;
    assign coff[1103] = 64'hffffcb75ffff8b48;
    assign coff[1104] = 64'hffffcb69ffff8b4d;
    assign coff[1105] = 64'hffffcb5effff8b52;
    assign coff[1106] = 64'hffffcb53ffff8b58;
    assign coff[1107] = 64'hffffcb47ffff8b5d;
    assign coff[1108] = 64'hffffcb3cffff8b62;
    assign coff[1109] = 64'hffffcb30ffff8b67;
    assign coff[1110] = 64'hffffcb25ffff8b6c;
    assign coff[1111] = 64'hffffcb19ffff8b71;
    assign coff[1112] = 64'hffffcb0effff8b77;
    assign coff[1113] = 64'hffffcb02ffff8b7c;
    assign coff[1114] = 64'hffffcaf7ffff8b81;
    assign coff[1115] = 64'hffffcaecffff8b86;
    assign coff[1116] = 64'hffffcae0ffff8b8b;
    assign coff[1117] = 64'hffffcad5ffff8b91;
    assign coff[1118] = 64'hffffcac9ffff8b96;
    assign coff[1119] = 64'hffffcabeffff8b9b;
    assign coff[1120] = 64'hffffcab2ffff8ba0;
    assign coff[1121] = 64'hffffcaa7ffff8ba6;
    assign coff[1122] = 64'hffffca9cffff8bab;
    assign coff[1123] = 64'hffffca90ffff8bb0;
    assign coff[1124] = 64'hffffca85ffff8bb5;
    assign coff[1125] = 64'hffffca79ffff8bbb;
    assign coff[1126] = 64'hffffca6effff8bc0;
    assign coff[1127] = 64'hffffca63ffff8bc5;
    assign coff[1128] = 64'hffffca57ffff8bca;
    assign coff[1129] = 64'hffffca4cffff8bd0;
    assign coff[1130] = 64'hffffca40ffff8bd5;
    assign coff[1131] = 64'hffffca35ffff8bda;
    assign coff[1132] = 64'hffffca29ffff8bdf;
    assign coff[1133] = 64'hffffca1effff8be5;
    assign coff[1134] = 64'hffffca13ffff8bea;
    assign coff[1135] = 64'hffffca07ffff8bef;
    assign coff[1136] = 64'hffffc9fcffff8bf5;
    assign coff[1137] = 64'hffffc9f1ffff8bfa;
    assign coff[1138] = 64'hffffc9e5ffff8bff;
    assign coff[1139] = 64'hffffc9daffff8c05;
    assign coff[1140] = 64'hffffc9ceffff8c0a;
    assign coff[1141] = 64'hffffc9c3ffff8c0f;
    assign coff[1142] = 64'hffffc9b8ffff8c15;
    assign coff[1143] = 64'hffffc9acffff8c1a;
    assign coff[1144] = 64'hffffc9a1ffff8c1f;
    assign coff[1145] = 64'hffffc995ffff8c25;
    assign coff[1146] = 64'hffffc98affff8c2a;
    assign coff[1147] = 64'hffffc97fffff8c2f;
    assign coff[1148] = 64'hffffc973ffff8c35;
    assign coff[1149] = 64'hffffc968ffff8c3a;
    assign coff[1150] = 64'hffffc95dffff8c3f;
    assign coff[1151] = 64'hffffc951ffff8c45;
    assign coff[1152] = 64'hffffc946ffff8c4a;
    assign coff[1153] = 64'hffffc93bffff8c4f;
    assign coff[1154] = 64'hffffc92fffff8c55;
    assign coff[1155] = 64'hffffc924ffff8c5a;
    assign coff[1156] = 64'hffffc918ffff8c60;
    assign coff[1157] = 64'hffffc90dffff8c65;
    assign coff[1158] = 64'hffffc902ffff8c6a;
    assign coff[1159] = 64'hffffc8f6ffff8c70;
    assign coff[1160] = 64'hffffc8ebffff8c75;
    assign coff[1161] = 64'hffffc8e0ffff8c7b;
    assign coff[1162] = 64'hffffc8d4ffff8c80;
    assign coff[1163] = 64'hffffc8c9ffff8c85;
    assign coff[1164] = 64'hffffc8beffff8c8b;
    assign coff[1165] = 64'hffffc8b2ffff8c90;
    assign coff[1166] = 64'hffffc8a7ffff8c96;
    assign coff[1167] = 64'hffffc89cffff8c9b;
    assign coff[1168] = 64'hffffc890ffff8ca1;
    assign coff[1169] = 64'hffffc885ffff8ca6;
    assign coff[1170] = 64'hffffc87affff8cab;
    assign coff[1171] = 64'hffffc86effff8cb1;
    assign coff[1172] = 64'hffffc863ffff8cb6;
    assign coff[1173] = 64'hffffc858ffff8cbc;
    assign coff[1174] = 64'hffffc84cffff8cc1;
    assign coff[1175] = 64'hffffc841ffff8cc7;
    assign coff[1176] = 64'hffffc836ffff8ccc;
    assign coff[1177] = 64'hffffc82bffff8cd2;
    assign coff[1178] = 64'hffffc81fffff8cd7;
    assign coff[1179] = 64'hffffc814ffff8cdd;
    assign coff[1180] = 64'hffffc809ffff8ce2;
    assign coff[1181] = 64'hffffc7fdffff8ce8;
    assign coff[1182] = 64'hffffc7f2ffff8ced;
    assign coff[1183] = 64'hffffc7e7ffff8cf3;
    assign coff[1184] = 64'hffffc7dbffff8cf8;
    assign coff[1185] = 64'hffffc7d0ffff8cfe;
    assign coff[1186] = 64'hffffc7c5ffff8d03;
    assign coff[1187] = 64'hffffc7baffff8d09;
    assign coff[1188] = 64'hffffc7aeffff8d0e;
    assign coff[1189] = 64'hffffc7a3ffff8d14;
    assign coff[1190] = 64'hffffc798ffff8d19;
    assign coff[1191] = 64'hffffc78cffff8d1f;
    assign coff[1192] = 64'hffffc781ffff8d24;
    assign coff[1193] = 64'hffffc776ffff8d2a;
    assign coff[1194] = 64'hffffc76bffff8d30;
    assign coff[1195] = 64'hffffc75fffff8d35;
    assign coff[1196] = 64'hffffc754ffff8d3b;
    assign coff[1197] = 64'hffffc749ffff8d40;
    assign coff[1198] = 64'hffffc73effff8d46;
    assign coff[1199] = 64'hffffc732ffff8d4b;
    assign coff[1200] = 64'hffffc727ffff8d51;
    assign coff[1201] = 64'hffffc71cffff8d57;
    assign coff[1202] = 64'hffffc710ffff8d5c;
    assign coff[1203] = 64'hffffc705ffff8d62;
    assign coff[1204] = 64'hffffc6faffff8d67;
    assign coff[1205] = 64'hffffc6efffff8d6d;
    assign coff[1206] = 64'hffffc6e3ffff8d73;
    assign coff[1207] = 64'hffffc6d8ffff8d78;
    assign coff[1208] = 64'hffffc6cdffff8d7e;
    assign coff[1209] = 64'hffffc6c2ffff8d83;
    assign coff[1210] = 64'hffffc6b7ffff8d89;
    assign coff[1211] = 64'hffffc6abffff8d8f;
    assign coff[1212] = 64'hffffc6a0ffff8d94;
    assign coff[1213] = 64'hffffc695ffff8d9a;
    assign coff[1214] = 64'hffffc68affff8da0;
    assign coff[1215] = 64'hffffc67effff8da5;
    assign coff[1216] = 64'hffffc673ffff8dab;
    assign coff[1217] = 64'hffffc668ffff8db0;
    assign coff[1218] = 64'hffffc65dffff8db6;
    assign coff[1219] = 64'hffffc651ffff8dbc;
    assign coff[1220] = 64'hffffc646ffff8dc1;
    assign coff[1221] = 64'hffffc63bffff8dc7;
    assign coff[1222] = 64'hffffc630ffff8dcd;
    assign coff[1223] = 64'hffffc625ffff8dd2;
    assign coff[1224] = 64'hffffc619ffff8dd8;
    assign coff[1225] = 64'hffffc60effff8dde;
    assign coff[1226] = 64'hffffc603ffff8de4;
    assign coff[1227] = 64'hffffc5f8ffff8de9;
    assign coff[1228] = 64'hffffc5edffff8def;
    assign coff[1229] = 64'hffffc5e1ffff8df5;
    assign coff[1230] = 64'hffffc5d6ffff8dfa;
    assign coff[1231] = 64'hffffc5cbffff8e00;
    assign coff[1232] = 64'hffffc5c0ffff8e06;
    assign coff[1233] = 64'hffffc5b5ffff8e0b;
    assign coff[1234] = 64'hffffc5a9ffff8e11;
    assign coff[1235] = 64'hffffc59effff8e17;
    assign coff[1236] = 64'hffffc593ffff8e1d;
    assign coff[1237] = 64'hffffc588ffff8e22;
    assign coff[1238] = 64'hffffc57dffff8e28;
    assign coff[1239] = 64'hffffc572ffff8e2e;
    assign coff[1240] = 64'hffffc566ffff8e34;
    assign coff[1241] = 64'hffffc55bffff8e39;
    assign coff[1242] = 64'hffffc550ffff8e3f;
    assign coff[1243] = 64'hffffc545ffff8e45;
    assign coff[1244] = 64'hffffc53affff8e4b;
    assign coff[1245] = 64'hffffc52fffff8e50;
    assign coff[1246] = 64'hffffc523ffff8e56;
    assign coff[1247] = 64'hffffc518ffff8e5c;
    assign coff[1248] = 64'hffffc50dffff8e62;
    assign coff[1249] = 64'hffffc502ffff8e68;
    assign coff[1250] = 64'hffffc4f7ffff8e6d;
    assign coff[1251] = 64'hffffc4ecffff8e73;
    assign coff[1252] = 64'hffffc4e0ffff8e79;
    assign coff[1253] = 64'hffffc4d5ffff8e7f;
    assign coff[1254] = 64'hffffc4caffff8e85;
    assign coff[1255] = 64'hffffc4bfffff8e8a;
    assign coff[1256] = 64'hffffc4b4ffff8e90;
    assign coff[1257] = 64'hffffc4a9ffff8e96;
    assign coff[1258] = 64'hffffc49effff8e9c;
    assign coff[1259] = 64'hffffc493ffff8ea2;
    assign coff[1260] = 64'hffffc487ffff8ea8;
    assign coff[1261] = 64'hffffc47cffff8ead;
    assign coff[1262] = 64'hffffc471ffff8eb3;
    assign coff[1263] = 64'hffffc466ffff8eb9;
    assign coff[1264] = 64'hffffc45bffff8ebf;
    assign coff[1265] = 64'hffffc450ffff8ec5;
    assign coff[1266] = 64'hffffc445ffff8ecb;
    assign coff[1267] = 64'hffffc43affff8ed1;
    assign coff[1268] = 64'hffffc42effff8ed6;
    assign coff[1269] = 64'hffffc423ffff8edc;
    assign coff[1270] = 64'hffffc418ffff8ee2;
    assign coff[1271] = 64'hffffc40dffff8ee8;
    assign coff[1272] = 64'hffffc402ffff8eee;
    assign coff[1273] = 64'hffffc3f7ffff8ef4;
    assign coff[1274] = 64'hffffc3ecffff8efa;
    assign coff[1275] = 64'hffffc3e1ffff8f00;
    assign coff[1276] = 64'hffffc3d6ffff8f06;
    assign coff[1277] = 64'hffffc3cbffff8f0b;
    assign coff[1278] = 64'hffffc3bfffff8f11;
    assign coff[1279] = 64'hffffc3b4ffff8f17;
    assign coff[1280] = 64'hffffc3a9ffff8f1d;
    assign coff[1281] = 64'hffffc39effff8f23;
    assign coff[1282] = 64'hffffc393ffff8f29;
    assign coff[1283] = 64'hffffc388ffff8f2f;
    assign coff[1284] = 64'hffffc37dffff8f35;
    assign coff[1285] = 64'hffffc372ffff8f3b;
    assign coff[1286] = 64'hffffc367ffff8f41;
    assign coff[1287] = 64'hffffc35cffff8f47;
    assign coff[1288] = 64'hffffc351ffff8f4d;
    assign coff[1289] = 64'hffffc346ffff8f53;
    assign coff[1290] = 64'hffffc33bffff8f59;
    assign coff[1291] = 64'hffffc330ffff8f5f;
    assign coff[1292] = 64'hffffc324ffff8f65;
    assign coff[1293] = 64'hffffc319ffff8f6b;
    assign coff[1294] = 64'hffffc30effff8f71;
    assign coff[1295] = 64'hffffc303ffff8f77;
    assign coff[1296] = 64'hffffc2f8ffff8f7d;
    assign coff[1297] = 64'hffffc2edffff8f83;
    assign coff[1298] = 64'hffffc2e2ffff8f89;
    assign coff[1299] = 64'hffffc2d7ffff8f8f;
    assign coff[1300] = 64'hffffc2ccffff8f95;
    assign coff[1301] = 64'hffffc2c1ffff8f9b;
    assign coff[1302] = 64'hffffc2b6ffff8fa1;
    assign coff[1303] = 64'hffffc2abffff8fa7;
    assign coff[1304] = 64'hffffc2a0ffff8fad;
    assign coff[1305] = 64'hffffc295ffff8fb3;
    assign coff[1306] = 64'hffffc28affff8fb9;
    assign coff[1307] = 64'hffffc27fffff8fbf;
    assign coff[1308] = 64'hffffc274ffff8fc5;
    assign coff[1309] = 64'hffffc269ffff8fcb;
    assign coff[1310] = 64'hffffc25effff8fd1;
    assign coff[1311] = 64'hffffc253ffff8fd7;
    assign coff[1312] = 64'hffffc248ffff8fdd;
    assign coff[1313] = 64'hffffc23dffff8fe3;
    assign coff[1314] = 64'hffffc232ffff8fe9;
    assign coff[1315] = 64'hffffc227ffff8fef;
    assign coff[1316] = 64'hffffc21cffff8ff5;
    assign coff[1317] = 64'hffffc211ffff8ffb;
    assign coff[1318] = 64'hffffc206ffff9001;
    assign coff[1319] = 64'hffffc1fbffff9007;
    assign coff[1320] = 64'hffffc1f0ffff900e;
    assign coff[1321] = 64'hffffc1e5ffff9014;
    assign coff[1322] = 64'hffffc1daffff901a;
    assign coff[1323] = 64'hffffc1cfffff9020;
    assign coff[1324] = 64'hffffc1c4ffff9026;
    assign coff[1325] = 64'hffffc1b9ffff902c;
    assign coff[1326] = 64'hffffc1aeffff9032;
    assign coff[1327] = 64'hffffc1a3ffff9038;
    assign coff[1328] = 64'hffffc198ffff903e;
    assign coff[1329] = 64'hffffc18dffff9045;
    assign coff[1330] = 64'hffffc182ffff904b;
    assign coff[1331] = 64'hffffc177ffff9051;
    assign coff[1332] = 64'hffffc16cffff9057;
    assign coff[1333] = 64'hffffc161ffff905d;
    assign coff[1334] = 64'hffffc156ffff9063;
    assign coff[1335] = 64'hffffc14bffff9069;
    assign coff[1336] = 64'hffffc140ffff9070;
    assign coff[1337] = 64'hffffc135ffff9076;
    assign coff[1338] = 64'hffffc12affff907c;
    assign coff[1339] = 64'hffffc11fffff9082;
    assign coff[1340] = 64'hffffc114ffff9088;
    assign coff[1341] = 64'hffffc10affff908e;
    assign coff[1342] = 64'hffffc0ffffff9095;
    assign coff[1343] = 64'hffffc0f4ffff909b;
    assign coff[1344] = 64'hffffc0e9ffff90a1;
    assign coff[1345] = 64'hffffc0deffff90a7;
    assign coff[1346] = 64'hffffc0d3ffff90ad;
    assign coff[1347] = 64'hffffc0c8ffff90b4;
    assign coff[1348] = 64'hffffc0bdffff90ba;
    assign coff[1349] = 64'hffffc0b2ffff90c0;
    assign coff[1350] = 64'hffffc0a7ffff90c6;
    assign coff[1351] = 64'hffffc09cffff90cc;
    assign coff[1352] = 64'hffffc091ffff90d3;
    assign coff[1353] = 64'hffffc086ffff90d9;
    assign coff[1354] = 64'hffffc07bffff90df;
    assign coff[1355] = 64'hffffc071ffff90e5;
    assign coff[1356] = 64'hffffc066ffff90ec;
    assign coff[1357] = 64'hffffc05bffff90f2;
    assign coff[1358] = 64'hffffc050ffff90f8;
    assign coff[1359] = 64'hffffc045ffff90fe;
    assign coff[1360] = 64'hffffc03affff9105;
    assign coff[1361] = 64'hffffc02fffff910b;
    assign coff[1362] = 64'hffffc024ffff9111;
    assign coff[1363] = 64'hffffc019ffff9117;
    assign coff[1364] = 64'hffffc00fffff911e;
    assign coff[1365] = 64'hffffc004ffff9124;
    assign coff[1366] = 64'hffffbff9ffff912a;
    assign coff[1367] = 64'hffffbfeeffff9131;
    assign coff[1368] = 64'hffffbfe3ffff9137;
    assign coff[1369] = 64'hffffbfd8ffff913d;
    assign coff[1370] = 64'hffffbfcdffff9143;
    assign coff[1371] = 64'hffffbfc2ffff914a;
    assign coff[1372] = 64'hffffbfb8ffff9150;
    assign coff[1373] = 64'hffffbfadffff9156;
    assign coff[1374] = 64'hffffbfa2ffff915d;
    assign coff[1375] = 64'hffffbf97ffff9163;
    assign coff[1376] = 64'hffffbf8cffff9169;
    assign coff[1377] = 64'hffffbf81ffff9170;
    assign coff[1378] = 64'hffffbf76ffff9176;
    assign coff[1379] = 64'hffffbf6bffff917c;
    assign coff[1380] = 64'hffffbf61ffff9183;
    assign coff[1381] = 64'hffffbf56ffff9189;
    assign coff[1382] = 64'hffffbf4bffff918f;
    assign coff[1383] = 64'hffffbf40ffff9196;
    assign coff[1384] = 64'hffffbf35ffff919c;
    assign coff[1385] = 64'hffffbf2affff91a2;
    assign coff[1386] = 64'hffffbf20ffff91a9;
    assign coff[1387] = 64'hffffbf15ffff91af;
    assign coff[1388] = 64'hffffbf0affff91b6;
    assign coff[1389] = 64'hffffbeffffff91bc;
    assign coff[1390] = 64'hffffbef4ffff91c2;
    assign coff[1391] = 64'hffffbee9ffff91c9;
    assign coff[1392] = 64'hffffbedfffff91cf;
    assign coff[1393] = 64'hffffbed4ffff91d6;
    assign coff[1394] = 64'hffffbec9ffff91dc;
    assign coff[1395] = 64'hffffbebeffff91e2;
    assign coff[1396] = 64'hffffbeb3ffff91e9;
    assign coff[1397] = 64'hffffbea9ffff91ef;
    assign coff[1398] = 64'hffffbe9effff91f6;
    assign coff[1399] = 64'hffffbe93ffff91fc;
    assign coff[1400] = 64'hffffbe88ffff9202;
    assign coff[1401] = 64'hffffbe7dffff9209;
    assign coff[1402] = 64'hffffbe73ffff920f;
    assign coff[1403] = 64'hffffbe68ffff9216;
    assign coff[1404] = 64'hffffbe5dffff921c;
    assign coff[1405] = 64'hffffbe52ffff9223;
    assign coff[1406] = 64'hffffbe47ffff9229;
    assign coff[1407] = 64'hffffbe3dffff922f;
    assign coff[1408] = 64'hffffbe32ffff9236;
    assign coff[1409] = 64'hffffbe27ffff923c;
    assign coff[1410] = 64'hffffbe1cffff9243;
    assign coff[1411] = 64'hffffbe12ffff9249;
    assign coff[1412] = 64'hffffbe07ffff9250;
    assign coff[1413] = 64'hffffbdfcffff9256;
    assign coff[1414] = 64'hffffbdf1ffff925d;
    assign coff[1415] = 64'hffffbde6ffff9263;
    assign coff[1416] = 64'hffffbddcffff926a;
    assign coff[1417] = 64'hffffbdd1ffff9270;
    assign coff[1418] = 64'hffffbdc6ffff9277;
    assign coff[1419] = 64'hffffbdbbffff927d;
    assign coff[1420] = 64'hffffbdb1ffff9284;
    assign coff[1421] = 64'hffffbda6ffff928a;
    assign coff[1422] = 64'hffffbd9bffff9291;
    assign coff[1423] = 64'hffffbd90ffff9297;
    assign coff[1424] = 64'hffffbd86ffff929e;
    assign coff[1425] = 64'hffffbd7bffff92a4;
    assign coff[1426] = 64'hffffbd70ffff92ab;
    assign coff[1427] = 64'hffffbd66ffff92b1;
    assign coff[1428] = 64'hffffbd5bffff92b8;
    assign coff[1429] = 64'hffffbd50ffff92bf;
    assign coff[1430] = 64'hffffbd45ffff92c5;
    assign coff[1431] = 64'hffffbd3bffff92cc;
    assign coff[1432] = 64'hffffbd30ffff92d2;
    assign coff[1433] = 64'hffffbd25ffff92d9;
    assign coff[1434] = 64'hffffbd1affff92df;
    assign coff[1435] = 64'hffffbd10ffff92e6;
    assign coff[1436] = 64'hffffbd05ffff92ec;
    assign coff[1437] = 64'hffffbcfaffff92f3;
    assign coff[1438] = 64'hffffbcf0ffff92fa;
    assign coff[1439] = 64'hffffbce5ffff9300;
    assign coff[1440] = 64'hffffbcdaffff9307;
    assign coff[1441] = 64'hffffbcd0ffff930d;
    assign coff[1442] = 64'hffffbcc5ffff9314;
    assign coff[1443] = 64'hffffbcbaffff931b;
    assign coff[1444] = 64'hffffbcafffff9321;
    assign coff[1445] = 64'hffffbca5ffff9328;
    assign coff[1446] = 64'hffffbc9affff932e;
    assign coff[1447] = 64'hffffbc8fffff9335;
    assign coff[1448] = 64'hffffbc85ffff933c;
    assign coff[1449] = 64'hffffbc7affff9342;
    assign coff[1450] = 64'hffffbc6fffff9349;
    assign coff[1451] = 64'hffffbc65ffff9350;
    assign coff[1452] = 64'hffffbc5affff9356;
    assign coff[1453] = 64'hffffbc4fffff935d;
    assign coff[1454] = 64'hffffbc45ffff9363;
    assign coff[1455] = 64'hffffbc3affff936a;
    assign coff[1456] = 64'hffffbc2fffff9371;
    assign coff[1457] = 64'hffffbc25ffff9377;
    assign coff[1458] = 64'hffffbc1affff937e;
    assign coff[1459] = 64'hffffbc0fffff9385;
    assign coff[1460] = 64'hffffbc05ffff938b;
    assign coff[1461] = 64'hffffbbfaffff9392;
    assign coff[1462] = 64'hffffbbefffff9399;
    assign coff[1463] = 64'hffffbbe5ffff939f;
    assign coff[1464] = 64'hffffbbdaffff93a6;
    assign coff[1465] = 64'hffffbbd0ffff93ad;
    assign coff[1466] = 64'hffffbbc5ffff93b4;
    assign coff[1467] = 64'hffffbbbaffff93ba;
    assign coff[1468] = 64'hffffbbb0ffff93c1;
    assign coff[1469] = 64'hffffbba5ffff93c8;
    assign coff[1470] = 64'hffffbb9affff93ce;
    assign coff[1471] = 64'hffffbb90ffff93d5;
    assign coff[1472] = 64'hffffbb85ffff93dc;
    assign coff[1473] = 64'hffffbb7bffff93e3;
    assign coff[1474] = 64'hffffbb70ffff93e9;
    assign coff[1475] = 64'hffffbb65ffff93f0;
    assign coff[1476] = 64'hffffbb5bffff93f7;
    assign coff[1477] = 64'hffffbb50ffff93fe;
    assign coff[1478] = 64'hffffbb46ffff9404;
    assign coff[1479] = 64'hffffbb3bffff940b;
    assign coff[1480] = 64'hffffbb30ffff9412;
    assign coff[1481] = 64'hffffbb26ffff9419;
    assign coff[1482] = 64'hffffbb1bffff941f;
    assign coff[1483] = 64'hffffbb11ffff9426;
    assign coff[1484] = 64'hffffbb06ffff942d;
    assign coff[1485] = 64'hffffbafbffff9434;
    assign coff[1486] = 64'hffffbaf1ffff943a;
    assign coff[1487] = 64'hffffbae6ffff9441;
    assign coff[1488] = 64'hffffbadcffff9448;
    assign coff[1489] = 64'hffffbad1ffff944f;
    assign coff[1490] = 64'hffffbac7ffff9456;
    assign coff[1491] = 64'hffffbabcffff945c;
    assign coff[1492] = 64'hffffbab1ffff9463;
    assign coff[1493] = 64'hffffbaa7ffff946a;
    assign coff[1494] = 64'hffffba9cffff9471;
    assign coff[1495] = 64'hffffba92ffff9478;
    assign coff[1496] = 64'hffffba87ffff947e;
    assign coff[1497] = 64'hffffba7dffff9485;
    assign coff[1498] = 64'hffffba72ffff948c;
    assign coff[1499] = 64'hffffba67ffff9493;
    assign coff[1500] = 64'hffffba5dffff949a;
    assign coff[1501] = 64'hffffba52ffff94a1;
    assign coff[1502] = 64'hffffba48ffff94a7;
    assign coff[1503] = 64'hffffba3dffff94ae;
    assign coff[1504] = 64'hffffba33ffff94b5;
    assign coff[1505] = 64'hffffba28ffff94bc;
    assign coff[1506] = 64'hffffba1effff94c3;
    assign coff[1507] = 64'hffffba13ffff94ca;
    assign coff[1508] = 64'hffffba09ffff94d0;
    assign coff[1509] = 64'hffffb9feffff94d7;
    assign coff[1510] = 64'hffffb9f4ffff94de;
    assign coff[1511] = 64'hffffb9e9ffff94e5;
    assign coff[1512] = 64'hffffb9dfffff94ec;
    assign coff[1513] = 64'hffffb9d4ffff94f3;
    assign coff[1514] = 64'hffffb9caffff94fa;
    assign coff[1515] = 64'hffffb9bfffff9501;
    assign coff[1516] = 64'hffffb9b5ffff9508;
    assign coff[1517] = 64'hffffb9aaffff950e;
    assign coff[1518] = 64'hffffb9a0ffff9515;
    assign coff[1519] = 64'hffffb995ffff951c;
    assign coff[1520] = 64'hffffb98bffff9523;
    assign coff[1521] = 64'hffffb980ffff952a;
    assign coff[1522] = 64'hffffb976ffff9531;
    assign coff[1523] = 64'hffffb96bffff9538;
    assign coff[1524] = 64'hffffb961ffff953f;
    assign coff[1525] = 64'hffffb956ffff9546;
    assign coff[1526] = 64'hffffb94cffff954d;
    assign coff[1527] = 64'hffffb941ffff9554;
    assign coff[1528] = 64'hffffb937ffff955b;
    assign coff[1529] = 64'hffffb92cffff9562;
    assign coff[1530] = 64'hffffb922ffff9569;
    assign coff[1531] = 64'hffffb917ffff9570;
    assign coff[1532] = 64'hffffb90dffff9577;
    assign coff[1533] = 64'hffffb902ffff957d;
    assign coff[1534] = 64'hffffb8f8ffff9584;
    assign coff[1535] = 64'hffffb8eeffff958b;
    assign coff[1536] = 64'hffffb8e3ffff9592;
    assign coff[1537] = 64'hffffb8d9ffff9599;
    assign coff[1538] = 64'hffffb8ceffff95a0;
    assign coff[1539] = 64'hffffb8c4ffff95a7;
    assign coff[1540] = 64'hffffb8b9ffff95ae;
    assign coff[1541] = 64'hffffb8afffff95b5;
    assign coff[1542] = 64'hffffb8a4ffff95bc;
    assign coff[1543] = 64'hffffb89affff95c3;
    assign coff[1544] = 64'hffffb890ffff95ca;
    assign coff[1545] = 64'hffffb885ffff95d1;
    assign coff[1546] = 64'hffffb87bffff95d8;
    assign coff[1547] = 64'hffffb870ffff95df;
    assign coff[1548] = 64'hffffb866ffff95e6;
    assign coff[1549] = 64'hffffb85bffff95ee;
    assign coff[1550] = 64'hffffb851ffff95f5;
    assign coff[1551] = 64'hffffb847ffff95fc;
    assign coff[1552] = 64'hffffb83cffff9603;
    assign coff[1553] = 64'hffffb832ffff960a;
    assign coff[1554] = 64'hffffb827ffff9611;
    assign coff[1555] = 64'hffffb81dffff9618;
    assign coff[1556] = 64'hffffb813ffff961f;
    assign coff[1557] = 64'hffffb808ffff9626;
    assign coff[1558] = 64'hffffb7feffff962d;
    assign coff[1559] = 64'hffffb7f3ffff9634;
    assign coff[1560] = 64'hffffb7e9ffff963b;
    assign coff[1561] = 64'hffffb7dfffff9642;
    assign coff[1562] = 64'hffffb7d4ffff9649;
    assign coff[1563] = 64'hffffb7caffff9650;
    assign coff[1564] = 64'hffffb7c0ffff9657;
    assign coff[1565] = 64'hffffb7b5ffff965f;
    assign coff[1566] = 64'hffffb7abffff9666;
    assign coff[1567] = 64'hffffb7a0ffff966d;
    assign coff[1568] = 64'hffffb796ffff9674;
    assign coff[1569] = 64'hffffb78cffff967b;
    assign coff[1570] = 64'hffffb781ffff9682;
    assign coff[1571] = 64'hffffb777ffff9689;
    assign coff[1572] = 64'hffffb76dffff9690;
    assign coff[1573] = 64'hffffb762ffff9697;
    assign coff[1574] = 64'hffffb758ffff969f;
    assign coff[1575] = 64'hffffb74effff96a6;
    assign coff[1576] = 64'hffffb743ffff96ad;
    assign coff[1577] = 64'hffffb739ffff96b4;
    assign coff[1578] = 64'hffffb72fffff96bb;
    assign coff[1579] = 64'hffffb724ffff96c2;
    assign coff[1580] = 64'hffffb71affff96c9;
    assign coff[1581] = 64'hffffb710ffff96d1;
    assign coff[1582] = 64'hffffb705ffff96d8;
    assign coff[1583] = 64'hffffb6fbffff96df;
    assign coff[1584] = 64'hffffb6f1ffff96e6;
    assign coff[1585] = 64'hffffb6e6ffff96ed;
    assign coff[1586] = 64'hffffb6dcffff96f4;
    assign coff[1587] = 64'hffffb6d2ffff96fc;
    assign coff[1588] = 64'hffffb6c7ffff9703;
    assign coff[1589] = 64'hffffb6bdffff970a;
    assign coff[1590] = 64'hffffb6b3ffff9711;
    assign coff[1591] = 64'hffffb6a8ffff9718;
    assign coff[1592] = 64'hffffb69effff9720;
    assign coff[1593] = 64'hffffb694ffff9727;
    assign coff[1594] = 64'hffffb68affff972e;
    assign coff[1595] = 64'hffffb67fffff9735;
    assign coff[1596] = 64'hffffb675ffff973c;
    assign coff[1597] = 64'hffffb66bffff9744;
    assign coff[1598] = 64'hffffb660ffff974b;
    assign coff[1599] = 64'hffffb656ffff9752;
    assign coff[1600] = 64'hffffb64cffff9759;
    assign coff[1601] = 64'hffffb642ffff9761;
    assign coff[1602] = 64'hffffb637ffff9768;
    assign coff[1603] = 64'hffffb62dffff976f;
    assign coff[1604] = 64'hffffb623ffff9776;
    assign coff[1605] = 64'hffffb619ffff977e;
    assign coff[1606] = 64'hffffb60effff9785;
    assign coff[1607] = 64'hffffb604ffff978c;
    assign coff[1608] = 64'hffffb5faffff9793;
    assign coff[1609] = 64'hffffb5f0ffff979b;
    assign coff[1610] = 64'hffffb5e5ffff97a2;
    assign coff[1611] = 64'hffffb5dbffff97a9;
    assign coff[1612] = 64'hffffb5d1ffff97b0;
    assign coff[1613] = 64'hffffb5c7ffff97b8;
    assign coff[1614] = 64'hffffb5bcffff97bf;
    assign coff[1615] = 64'hffffb5b2ffff97c6;
    assign coff[1616] = 64'hffffb5a8ffff97ce;
    assign coff[1617] = 64'hffffb59effff97d5;
    assign coff[1618] = 64'hffffb593ffff97dc;
    assign coff[1619] = 64'hffffb589ffff97e4;
    assign coff[1620] = 64'hffffb57fffff97eb;
    assign coff[1621] = 64'hffffb575ffff97f2;
    assign coff[1622] = 64'hffffb56bffff97fa;
    assign coff[1623] = 64'hffffb560ffff9801;
    assign coff[1624] = 64'hffffb556ffff9808;
    assign coff[1625] = 64'hffffb54cffff9810;
    assign coff[1626] = 64'hffffb542ffff9817;
    assign coff[1627] = 64'hffffb538ffff981e;
    assign coff[1628] = 64'hffffb52dffff9826;
    assign coff[1629] = 64'hffffb523ffff982d;
    assign coff[1630] = 64'hffffb519ffff9834;
    assign coff[1631] = 64'hffffb50fffff983c;
    assign coff[1632] = 64'hffffb505ffff9843;
    assign coff[1633] = 64'hffffb4faffff984a;
    assign coff[1634] = 64'hffffb4f0ffff9852;
    assign coff[1635] = 64'hffffb4e6ffff9859;
    assign coff[1636] = 64'hffffb4dcffff9860;
    assign coff[1637] = 64'hffffb4d2ffff9868;
    assign coff[1638] = 64'hffffb4c8ffff986f;
    assign coff[1639] = 64'hffffb4bdffff9877;
    assign coff[1640] = 64'hffffb4b3ffff987e;
    assign coff[1641] = 64'hffffb4a9ffff9885;
    assign coff[1642] = 64'hffffb49fffff988d;
    assign coff[1643] = 64'hffffb495ffff9894;
    assign coff[1644] = 64'hffffb48bffff989c;
    assign coff[1645] = 64'hffffb480ffff98a3;
    assign coff[1646] = 64'hffffb476ffff98aa;
    assign coff[1647] = 64'hffffb46cffff98b2;
    assign coff[1648] = 64'hffffb462ffff98b9;
    assign coff[1649] = 64'hffffb458ffff98c1;
    assign coff[1650] = 64'hffffb44effff98c8;
    assign coff[1651] = 64'hffffb444ffff98d0;
    assign coff[1652] = 64'hffffb439ffff98d7;
    assign coff[1653] = 64'hffffb42fffff98de;
    assign coff[1654] = 64'hffffb425ffff98e6;
    assign coff[1655] = 64'hffffb41bffff98ed;
    assign coff[1656] = 64'hffffb411ffff98f5;
    assign coff[1657] = 64'hffffb407ffff98fc;
    assign coff[1658] = 64'hffffb3fdffff9904;
    assign coff[1659] = 64'hffffb3f3ffff990b;
    assign coff[1660] = 64'hffffb3e9ffff9913;
    assign coff[1661] = 64'hffffb3deffff991a;
    assign coff[1662] = 64'hffffb3d4ffff9922;
    assign coff[1663] = 64'hffffb3caffff9929;
    assign coff[1664] = 64'hffffb3c0ffff9930;
    assign coff[1665] = 64'hffffb3b6ffff9938;
    assign coff[1666] = 64'hffffb3acffff993f;
    assign coff[1667] = 64'hffffb3a2ffff9947;
    assign coff[1668] = 64'hffffb398ffff994e;
    assign coff[1669] = 64'hffffb38effff9956;
    assign coff[1670] = 64'hffffb384ffff995d;
    assign coff[1671] = 64'hffffb37affff9965;
    assign coff[1672] = 64'hffffb36fffff996d;
    assign coff[1673] = 64'hffffb365ffff9974;
    assign coff[1674] = 64'hffffb35bffff997c;
    assign coff[1675] = 64'hffffb351ffff9983;
    assign coff[1676] = 64'hffffb347ffff998b;
    assign coff[1677] = 64'hffffb33dffff9992;
    assign coff[1678] = 64'hffffb333ffff999a;
    assign coff[1679] = 64'hffffb329ffff99a1;
    assign coff[1680] = 64'hffffb31fffff99a9;
    assign coff[1681] = 64'hffffb315ffff99b0;
    assign coff[1682] = 64'hffffb30bffff99b8;
    assign coff[1683] = 64'hffffb301ffff99bf;
    assign coff[1684] = 64'hffffb2f7ffff99c7;
    assign coff[1685] = 64'hffffb2edffff99cf;
    assign coff[1686] = 64'hffffb2e3ffff99d6;
    assign coff[1687] = 64'hffffb2d9ffff99de;
    assign coff[1688] = 64'hffffb2cfffff99e5;
    assign coff[1689] = 64'hffffb2c5ffff99ed;
    assign coff[1690] = 64'hffffb2bbffff99f4;
    assign coff[1691] = 64'hffffb2b1ffff99fc;
    assign coff[1692] = 64'hffffb2a7ffff9a04;
    assign coff[1693] = 64'hffffb29dffff9a0b;
    assign coff[1694] = 64'hffffb293ffff9a13;
    assign coff[1695] = 64'hffffb289ffff9a1a;
    assign coff[1696] = 64'hffffb27fffff9a22;
    assign coff[1697] = 64'hffffb275ffff9a2a;
    assign coff[1698] = 64'hffffb26bffff9a31;
    assign coff[1699] = 64'hffffb261ffff9a39;
    assign coff[1700] = 64'hffffb257ffff9a40;
    assign coff[1701] = 64'hffffb24dffff9a48;
    assign coff[1702] = 64'hffffb243ffff9a50;
    assign coff[1703] = 64'hffffb239ffff9a57;
    assign coff[1704] = 64'hffffb22fffff9a5f;
    assign coff[1705] = 64'hffffb225ffff9a67;
    assign coff[1706] = 64'hffffb21bffff9a6e;
    assign coff[1707] = 64'hffffb211ffff9a76;
    assign coff[1708] = 64'hffffb207ffff9a7e;
    assign coff[1709] = 64'hffffb1fdffff9a85;
    assign coff[1710] = 64'hffffb1f3ffff9a8d;
    assign coff[1711] = 64'hffffb1e9ffff9a95;
    assign coff[1712] = 64'hffffb1dfffff9a9c;
    assign coff[1713] = 64'hffffb1d5ffff9aa4;
    assign coff[1714] = 64'hffffb1cbffff9aac;
    assign coff[1715] = 64'hffffb1c1ffff9ab3;
    assign coff[1716] = 64'hffffb1b7ffff9abb;
    assign coff[1717] = 64'hffffb1adffff9ac3;
    assign coff[1718] = 64'hffffb1a3ffff9aca;
    assign coff[1719] = 64'hffffb199ffff9ad2;
    assign coff[1720] = 64'hffffb18fffff9ada;
    assign coff[1721] = 64'hffffb186ffff9ae1;
    assign coff[1722] = 64'hffffb17cffff9ae9;
    assign coff[1723] = 64'hffffb172ffff9af1;
    assign coff[1724] = 64'hffffb168ffff9af9;
    assign coff[1725] = 64'hffffb15effff9b00;
    assign coff[1726] = 64'hffffb154ffff9b08;
    assign coff[1727] = 64'hffffb14affff9b10;
    assign coff[1728] = 64'hffffb140ffff9b17;
    assign coff[1729] = 64'hffffb136ffff9b1f;
    assign coff[1730] = 64'hffffb12cffff9b27;
    assign coff[1731] = 64'hffffb122ffff9b2f;
    assign coff[1732] = 64'hffffb118ffff9b36;
    assign coff[1733] = 64'hffffb10fffff9b3e;
    assign coff[1734] = 64'hffffb105ffff9b46;
    assign coff[1735] = 64'hffffb0fbffff9b4e;
    assign coff[1736] = 64'hffffb0f1ffff9b55;
    assign coff[1737] = 64'hffffb0e7ffff9b5d;
    assign coff[1738] = 64'hffffb0ddffff9b65;
    assign coff[1739] = 64'hffffb0d3ffff9b6d;
    assign coff[1740] = 64'hffffb0c9ffff9b75;
    assign coff[1741] = 64'hffffb0c0ffff9b7c;
    assign coff[1742] = 64'hffffb0b6ffff9b84;
    assign coff[1743] = 64'hffffb0acffff9b8c;
    assign coff[1744] = 64'hffffb0a2ffff9b94;
    assign coff[1745] = 64'hffffb098ffff9b9b;
    assign coff[1746] = 64'hffffb08effff9ba3;
    assign coff[1747] = 64'hffffb084ffff9bab;
    assign coff[1748] = 64'hffffb07bffff9bb3;
    assign coff[1749] = 64'hffffb071ffff9bbb;
    assign coff[1750] = 64'hffffb067ffff9bc2;
    assign coff[1751] = 64'hffffb05dffff9bca;
    assign coff[1752] = 64'hffffb053ffff9bd2;
    assign coff[1753] = 64'hffffb049ffff9bda;
    assign coff[1754] = 64'hffffb040ffff9be2;
    assign coff[1755] = 64'hffffb036ffff9bea;
    assign coff[1756] = 64'hffffb02cffff9bf1;
    assign coff[1757] = 64'hffffb022ffff9bf9;
    assign coff[1758] = 64'hffffb018ffff9c01;
    assign coff[1759] = 64'hffffb00effff9c09;
    assign coff[1760] = 64'hffffb005ffff9c11;
    assign coff[1761] = 64'hffffaffbffff9c19;
    assign coff[1762] = 64'hffffaff1ffff9c21;
    assign coff[1763] = 64'hffffafe7ffff9c28;
    assign coff[1764] = 64'hffffafddffff9c30;
    assign coff[1765] = 64'hffffafd4ffff9c38;
    assign coff[1766] = 64'hffffafcaffff9c40;
    assign coff[1767] = 64'hffffafc0ffff9c48;
    assign coff[1768] = 64'hffffafb6ffff9c50;
    assign coff[1769] = 64'hffffafacffff9c58;
    assign coff[1770] = 64'hffffafa3ffff9c60;
    assign coff[1771] = 64'hffffaf99ffff9c67;
    assign coff[1772] = 64'hffffaf8fffff9c6f;
    assign coff[1773] = 64'hffffaf85ffff9c77;
    assign coff[1774] = 64'hffffaf7cffff9c7f;
    assign coff[1775] = 64'hffffaf72ffff9c87;
    assign coff[1776] = 64'hffffaf68ffff9c8f;
    assign coff[1777] = 64'hffffaf5effff9c97;
    assign coff[1778] = 64'hffffaf54ffff9c9f;
    assign coff[1779] = 64'hffffaf4bffff9ca7;
    assign coff[1780] = 64'hffffaf41ffff9caf;
    assign coff[1781] = 64'hffffaf37ffff9cb7;
    assign coff[1782] = 64'hffffaf2dffff9cbe;
    assign coff[1783] = 64'hffffaf24ffff9cc6;
    assign coff[1784] = 64'hffffaf1affff9cce;
    assign coff[1785] = 64'hffffaf10ffff9cd6;
    assign coff[1786] = 64'hffffaf07ffff9cde;
    assign coff[1787] = 64'hffffaefdffff9ce6;
    assign coff[1788] = 64'hffffaef3ffff9cee;
    assign coff[1789] = 64'hffffaee9ffff9cf6;
    assign coff[1790] = 64'hffffaee0ffff9cfe;
    assign coff[1791] = 64'hffffaed6ffff9d06;
    assign coff[1792] = 64'hffffaeccffff9d0e;
    assign coff[1793] = 64'hffffaec2ffff9d16;
    assign coff[1794] = 64'hffffaeb9ffff9d1e;
    assign coff[1795] = 64'hffffaeafffff9d26;
    assign coff[1796] = 64'hffffaea5ffff9d2e;
    assign coff[1797] = 64'hffffae9cffff9d36;
    assign coff[1798] = 64'hffffae92ffff9d3e;
    assign coff[1799] = 64'hffffae88ffff9d46;
    assign coff[1800] = 64'hffffae7fffff9d4e;
    assign coff[1801] = 64'hffffae75ffff9d56;
    assign coff[1802] = 64'hffffae6bffff9d5e;
    assign coff[1803] = 64'hffffae62ffff9d66;
    assign coff[1804] = 64'hffffae58ffff9d6e;
    assign coff[1805] = 64'hffffae4effff9d76;
    assign coff[1806] = 64'hffffae45ffff9d7e;
    assign coff[1807] = 64'hffffae3bffff9d86;
    assign coff[1808] = 64'hffffae31ffff9d8e;
    assign coff[1809] = 64'hffffae28ffff9d96;
    assign coff[1810] = 64'hffffae1effff9d9e;
    assign coff[1811] = 64'hffffae14ffff9da6;
    assign coff[1812] = 64'hffffae0bffff9dae;
    assign coff[1813] = 64'hffffae01ffff9db6;
    assign coff[1814] = 64'hffffadf7ffff9dbe;
    assign coff[1815] = 64'hffffadeeffff9dc6;
    assign coff[1816] = 64'hffffade4ffff9dce;
    assign coff[1817] = 64'hffffaddaffff9dd6;
    assign coff[1818] = 64'hffffadd1ffff9ddf;
    assign coff[1819] = 64'hffffadc7ffff9de7;
    assign coff[1820] = 64'hffffadbdffff9def;
    assign coff[1821] = 64'hffffadb4ffff9df7;
    assign coff[1822] = 64'hffffadaaffff9dff;
    assign coff[1823] = 64'hffffada1ffff9e07;
    assign coff[1824] = 64'hffffad97ffff9e0f;
    assign coff[1825] = 64'hffffad8dffff9e17;
    assign coff[1826] = 64'hffffad84ffff9e1f;
    assign coff[1827] = 64'hffffad7affff9e27;
    assign coff[1828] = 64'hffffad70ffff9e2f;
    assign coff[1829] = 64'hffffad67ffff9e37;
    assign coff[1830] = 64'hffffad5dffff9e40;
    assign coff[1831] = 64'hffffad54ffff9e48;
    assign coff[1832] = 64'hffffad4affff9e50;
    assign coff[1833] = 64'hffffad41ffff9e58;
    assign coff[1834] = 64'hffffad37ffff9e60;
    assign coff[1835] = 64'hffffad2dffff9e68;
    assign coff[1836] = 64'hffffad24ffff9e70;
    assign coff[1837] = 64'hffffad1affff9e78;
    assign coff[1838] = 64'hffffad11ffff9e81;
    assign coff[1839] = 64'hffffad07ffff9e89;
    assign coff[1840] = 64'hffffacfdffff9e91;
    assign coff[1841] = 64'hffffacf4ffff9e99;
    assign coff[1842] = 64'hffffaceaffff9ea1;
    assign coff[1843] = 64'hfffface1ffff9ea9;
    assign coff[1844] = 64'hffffacd7ffff9eb2;
    assign coff[1845] = 64'hffffacceffff9eba;
    assign coff[1846] = 64'hffffacc4ffff9ec2;
    assign coff[1847] = 64'hffffacbbffff9eca;
    assign coff[1848] = 64'hffffacb1ffff9ed2;
    assign coff[1849] = 64'hffffaca8ffff9eda;
    assign coff[1850] = 64'hffffac9effff9ee3;
    assign coff[1851] = 64'hffffac94ffff9eeb;
    assign coff[1852] = 64'hffffac8bffff9ef3;
    assign coff[1853] = 64'hffffac81ffff9efb;
    assign coff[1854] = 64'hffffac78ffff9f03;
    assign coff[1855] = 64'hffffac6effff9f0c;
    assign coff[1856] = 64'hffffac65ffff9f14;
    assign coff[1857] = 64'hffffac5bffff9f1c;
    assign coff[1858] = 64'hffffac52ffff9f24;
    assign coff[1859] = 64'hffffac48ffff9f2c;
    assign coff[1860] = 64'hffffac3fffff9f35;
    assign coff[1861] = 64'hffffac35ffff9f3d;
    assign coff[1862] = 64'hffffac2cffff9f45;
    assign coff[1863] = 64'hffffac22ffff9f4d;
    assign coff[1864] = 64'hffffac19ffff9f56;
    assign coff[1865] = 64'hffffac0fffff9f5e;
    assign coff[1866] = 64'hffffac06ffff9f66;
    assign coff[1867] = 64'hffffabfcffff9f6e;
    assign coff[1868] = 64'hffffabf3ffff9f77;
    assign coff[1869] = 64'hffffabe9ffff9f7f;
    assign coff[1870] = 64'hffffabe0ffff9f87;
    assign coff[1871] = 64'hffffabd6ffff9f8f;
    assign coff[1872] = 64'hffffabcdffff9f98;
    assign coff[1873] = 64'hffffabc4ffff9fa0;
    assign coff[1874] = 64'hffffabbaffff9fa8;
    assign coff[1875] = 64'hffffabb1ffff9fb0;
    assign coff[1876] = 64'hffffaba7ffff9fb9;
    assign coff[1877] = 64'hffffab9effff9fc1;
    assign coff[1878] = 64'hffffab94ffff9fc9;
    assign coff[1879] = 64'hffffab8bffff9fd2;
    assign coff[1880] = 64'hffffab81ffff9fda;
    assign coff[1881] = 64'hffffab78ffff9fe2;
    assign coff[1882] = 64'hffffab6fffff9fea;
    assign coff[1883] = 64'hffffab65ffff9ff3;
    assign coff[1884] = 64'hffffab5cffff9ffb;
    assign coff[1885] = 64'hffffab52ffffa003;
    assign coff[1886] = 64'hffffab49ffffa00c;
    assign coff[1887] = 64'hffffab3fffffa014;
    assign coff[1888] = 64'hffffab36ffffa01c;
    assign coff[1889] = 64'hffffab2dffffa025;
    assign coff[1890] = 64'hffffab23ffffa02d;
    assign coff[1891] = 64'hffffab1affffa035;
    assign coff[1892] = 64'hffffab10ffffa03e;
    assign coff[1893] = 64'hffffab07ffffa046;
    assign coff[1894] = 64'hffffaafeffffa04e;
    assign coff[1895] = 64'hffffaaf4ffffa057;
    assign coff[1896] = 64'hffffaaebffffa05f;
    assign coff[1897] = 64'hffffaae1ffffa067;
    assign coff[1898] = 64'hffffaad8ffffa070;
    assign coff[1899] = 64'hffffaacfffffa078;
    assign coff[1900] = 64'hffffaac5ffffa080;
    assign coff[1901] = 64'hffffaabcffffa089;
    assign coff[1902] = 64'hffffaab2ffffa091;
    assign coff[1903] = 64'hffffaaa9ffffa09a;
    assign coff[1904] = 64'hffffaaa0ffffa0a2;
    assign coff[1905] = 64'hffffaa96ffffa0aa;
    assign coff[1906] = 64'hffffaa8dffffa0b3;
    assign coff[1907] = 64'hffffaa84ffffa0bb;
    assign coff[1908] = 64'hffffaa7affffa0c4;
    assign coff[1909] = 64'hffffaa71ffffa0cc;
    assign coff[1910] = 64'hffffaa68ffffa0d4;
    assign coff[1911] = 64'hffffaa5effffa0dd;
    assign coff[1912] = 64'hffffaa55ffffa0e5;
    assign coff[1913] = 64'hffffaa4cffffa0ee;
    assign coff[1914] = 64'hffffaa42ffffa0f6;
    assign coff[1915] = 64'hffffaa39ffffa0fe;
    assign coff[1916] = 64'hffffaa30ffffa107;
    assign coff[1917] = 64'hffffaa26ffffa10f;
    assign coff[1918] = 64'hffffaa1dffffa118;
    assign coff[1919] = 64'hffffaa14ffffa120;
    assign coff[1920] = 64'hffffaa0affffa129;
    assign coff[1921] = 64'hffffaa01ffffa131;
    assign coff[1922] = 64'hffffa9f8ffffa139;
    assign coff[1923] = 64'hffffa9eeffffa142;
    assign coff[1924] = 64'hffffa9e5ffffa14a;
    assign coff[1925] = 64'hffffa9dcffffa153;
    assign coff[1926] = 64'hffffa9d3ffffa15b;
    assign coff[1927] = 64'hffffa9c9ffffa164;
    assign coff[1928] = 64'hffffa9c0ffffa16c;
    assign coff[1929] = 64'hffffa9b7ffffa175;
    assign coff[1930] = 64'hffffa9adffffa17d;
    assign coff[1931] = 64'hffffa9a4ffffa186;
    assign coff[1932] = 64'hffffa99bffffa18e;
    assign coff[1933] = 64'hffffa992ffffa197;
    assign coff[1934] = 64'hffffa988ffffa19f;
    assign coff[1935] = 64'hffffa97fffffa1a8;
    assign coff[1936] = 64'hffffa976ffffa1b0;
    assign coff[1937] = 64'hffffa96dffffa1b8;
    assign coff[1938] = 64'hffffa963ffffa1c1;
    assign coff[1939] = 64'hffffa95affffa1c9;
    assign coff[1940] = 64'hffffa951ffffa1d2;
    assign coff[1941] = 64'hffffa948ffffa1db;
    assign coff[1942] = 64'hffffa93effffa1e3;
    assign coff[1943] = 64'hffffa935ffffa1ec;
    assign coff[1944] = 64'hffffa92cffffa1f4;
    assign coff[1945] = 64'hffffa923ffffa1fd;
    assign coff[1946] = 64'hffffa919ffffa205;
    assign coff[1947] = 64'hffffa910ffffa20e;
    assign coff[1948] = 64'hffffa907ffffa216;
    assign coff[1949] = 64'hffffa8feffffa21f;
    assign coff[1950] = 64'hffffa8f4ffffa227;
    assign coff[1951] = 64'hffffa8ebffffa230;
    assign coff[1952] = 64'hffffa8e2ffffa238;
    assign coff[1953] = 64'hffffa8d9ffffa241;
    assign coff[1954] = 64'hffffa8d0ffffa249;
    assign coff[1955] = 64'hffffa8c6ffffa252;
    assign coff[1956] = 64'hffffa8bdffffa25b;
    assign coff[1957] = 64'hffffa8b4ffffa263;
    assign coff[1958] = 64'hffffa8abffffa26c;
    assign coff[1959] = 64'hffffa8a2ffffa274;
    assign coff[1960] = 64'hffffa899ffffa27d;
    assign coff[1961] = 64'hffffa88fffffa286;
    assign coff[1962] = 64'hffffa886ffffa28e;
    assign coff[1963] = 64'hffffa87dffffa297;
    assign coff[1964] = 64'hffffa874ffffa29f;
    assign coff[1965] = 64'hffffa86bffffa2a8;
    assign coff[1966] = 64'hffffa861ffffa2b0;
    assign coff[1967] = 64'hffffa858ffffa2b9;
    assign coff[1968] = 64'hffffa84fffffa2c2;
    assign coff[1969] = 64'hffffa846ffffa2ca;
    assign coff[1970] = 64'hffffa83dffffa2d3;
    assign coff[1971] = 64'hffffa834ffffa2dc;
    assign coff[1972] = 64'hffffa82bffffa2e4;
    assign coff[1973] = 64'hffffa821ffffa2ed;
    assign coff[1974] = 64'hffffa818ffffa2f5;
    assign coff[1975] = 64'hffffa80fffffa2fe;
    assign coff[1976] = 64'hffffa806ffffa307;
    assign coff[1977] = 64'hffffa7fdffffa30f;
    assign coff[1978] = 64'hffffa7f4ffffa318;
    assign coff[1979] = 64'hffffa7ebffffa321;
    assign coff[1980] = 64'hffffa7e2ffffa329;
    assign coff[1981] = 64'hffffa7d8ffffa332;
    assign coff[1982] = 64'hffffa7cfffffa33b;
    assign coff[1983] = 64'hffffa7c6ffffa343;
    assign coff[1984] = 64'hffffa7bdffffa34c;
    assign coff[1985] = 64'hffffa7b4ffffa355;
    assign coff[1986] = 64'hffffa7abffffa35d;
    assign coff[1987] = 64'hffffa7a2ffffa366;
    assign coff[1988] = 64'hffffa799ffffa36f;
    assign coff[1989] = 64'hffffa790ffffa377;
    assign coff[1990] = 64'hffffa787ffffa380;
    assign coff[1991] = 64'hffffa77effffa389;
    assign coff[1992] = 64'hffffa774ffffa391;
    assign coff[1993] = 64'hffffa76bffffa39a;
    assign coff[1994] = 64'hffffa762ffffa3a3;
    assign coff[1995] = 64'hffffa759ffffa3ab;
    assign coff[1996] = 64'hffffa750ffffa3b4;
    assign coff[1997] = 64'hffffa747ffffa3bd;
    assign coff[1998] = 64'hffffa73effffa3c6;
    assign coff[1999] = 64'hffffa735ffffa3ce;
    assign coff[2000] = 64'hffffa72cffffa3d7;
    assign coff[2001] = 64'hffffa723ffffa3e0;
    assign coff[2002] = 64'hffffa71affffa3e8;
    assign coff[2003] = 64'hffffa711ffffa3f1;
    assign coff[2004] = 64'hffffa708ffffa3fa;
    assign coff[2005] = 64'hffffa6ffffffa403;
    assign coff[2006] = 64'hffffa6f6ffffa40b;
    assign coff[2007] = 64'hffffa6edffffa414;
    assign coff[2008] = 64'hffffa6e4ffffa41d;
    assign coff[2009] = 64'hffffa6dbffffa426;
    assign coff[2010] = 64'hffffa6d2ffffa42e;
    assign coff[2011] = 64'hffffa6c9ffffa437;
    assign coff[2012] = 64'hffffa6c0ffffa440;
    assign coff[2013] = 64'hffffa6b7ffffa449;
    assign coff[2014] = 64'hffffa6aeffffa451;
    assign coff[2015] = 64'hffffa6a5ffffa45a;
    assign coff[2016] = 64'hffffa69cffffa463;
    assign coff[2017] = 64'hffffa693ffffa46c;
    assign coff[2018] = 64'hffffa68affffa474;
    assign coff[2019] = 64'hffffa681ffffa47d;
    assign coff[2020] = 64'hffffa678ffffa486;
    assign coff[2021] = 64'hffffa66fffffa48f;
    assign coff[2022] = 64'hffffa666ffffa498;
    assign coff[2023] = 64'hffffa65dffffa4a0;
    assign coff[2024] = 64'hffffa654ffffa4a9;
    assign coff[2025] = 64'hffffa64bffffa4b2;
    assign coff[2026] = 64'hffffa642ffffa4bb;
    assign coff[2027] = 64'hffffa639ffffa4c4;
    assign coff[2028] = 64'hffffa630ffffa4cc;
    assign coff[2029] = 64'hffffa627ffffa4d5;
    assign coff[2030] = 64'hffffa61effffa4de;
    assign coff[2031] = 64'hffffa615ffffa4e7;
    assign coff[2032] = 64'hffffa60cffffa4f0;
    assign coff[2033] = 64'hffffa603ffffa4f9;
    assign coff[2034] = 64'hffffa5faffffa501;
    assign coff[2035] = 64'hffffa5f1ffffa50a;
    assign coff[2036] = 64'hffffa5e8ffffa513;
    assign coff[2037] = 64'hffffa5dfffffa51c;
    assign coff[2038] = 64'hffffa5d7ffffa525;
    assign coff[2039] = 64'hffffa5ceffffa52e;
    assign coff[2040] = 64'hffffa5c5ffffa537;
    assign coff[2041] = 64'hffffa5bcffffa53f;
    assign coff[2042] = 64'hffffa5b3ffffa548;
    assign coff[2043] = 64'hffffa5aaffffa551;
    assign coff[2044] = 64'hffffa5a1ffffa55a;
    assign coff[2045] = 64'hffffa598ffffa563;
    assign coff[2046] = 64'hffffa58fffffa56c;
    assign coff[2047] = 64'hffffa586ffffa575;




    always_ff @(posedge clk, negedge rst_n) begin
        if(~rst_n) begin
            data_o_col1 <= 'b0;
            data_o_col2 <= 'b0;
        end else begin
            if ((addr_col1 == 'd0 || addr_col1 == 'd1024) && (valid == 1)) begin
                data_o_col1 <= coff[addr_col1];
                data_o_col2 <= 'b0;
            end else if(valid == 1) begin
                data_o_col1 <= coff[addr_col1];
                data_o_col2 <= coff[addr_col2];
            end else begin
                data_o_col1 <= 'b0;
                data_o_col2 <= 'b0;
            end       
        end
    end


endmodule