`timescale 1ns/1ps
module rom_2
(
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic                     valid,
    input  logic [10:0]              addr_i,
    output logic [255:0]              data_o
);

    logic [255:0] coff[2047:0];

    assign coff[0   ] = 256'h00007fff00000000ffff80010000000000007fff00000000ffff800100000000;
    assign coff[1   ] = 256'h00000000ffff80010000000000007fff00000000ffff80010000000000007fff;
    assign coff[2   ] = 256'h00005a82ffffa57effffa57e00005a8200005a82ffffa57effffa57e00005a82;
    assign coff[3   ] = 256'hffffa57effffa57e00005a8200005a82ffffa57effffa57e00005a8200005a82;
    assign coff[4   ] = 256'h00007642ffffcf04ffff89be000030fc00007642ffffcf04ffff89be000030fc;
    assign coff[5   ] = 256'hffffcf04ffff89be000030fc00007642ffffcf04ffff89be000030fc00007642;
    assign coff[6   ] = 256'h000030fcffff89beffffcf0400007642000030fcffff89beffffcf0400007642;
    assign coff[7   ] = 256'hffff89beffffcf0400007642000030fcffff89beffffcf0400007642000030fc;
    assign coff[8   ] = 256'h00007d8affffe707ffff8276000018f900007d8affffe707ffff8276000018f9;
    assign coff[9   ] = 256'hffffe707ffff8276000018f900007d8affffe707ffff8276000018f900007d8a;
    assign coff[10  ] = 256'h0000471dffff9592ffffb8e300006a6e0000471dffff9592ffffb8e300006a6e;
    assign coff[11  ] = 256'hffff9592ffffb8e300006a6e0000471dffff9592ffffb8e300006a6e0000471d;
    assign coff[12  ] = 256'h00006a6effffb8e3ffff95920000471d00006a6effffb8e3ffff95920000471d;
    assign coff[13  ] = 256'hffffb8e3ffff95920000471d00006a6effffb8e3ffff95920000471d00006a6e;
    assign coff[14  ] = 256'h000018f9ffff8276ffffe70700007d8a000018f9ffff8276ffffe70700007d8a;
    assign coff[15  ] = 256'hffff8276ffffe70700007d8a000018f9ffff8276ffffe70700007d8a000018f9;
    assign coff[16  ] = 256'h00007f62fffff374ffff809e00000c8c00007f62fffff374ffff809e00000c8c;
    assign coff[17  ] = 256'hfffff374ffff809e00000c8c00007f62fffff374ffff809e00000c8c00007f62;
    assign coff[18  ] = 256'h00005134ffff9d0effffaecc000062f200005134ffff9d0effffaecc000062f2;
    assign coff[19  ] = 256'hffff9d0effffaecc000062f200005134ffff9d0effffaecc000062f200005134;
    assign coff[20  ] = 256'h000070e3ffffc3a9ffff8f1d00003c57000070e3ffffc3a9ffff8f1d00003c57;
    assign coff[21  ] = 256'hffffc3a9ffff8f1d00003c57000070e3ffffc3a9ffff8f1d00003c57000070e3;
    assign coff[22  ] = 256'h00002528ffff8583ffffdad800007a7d00002528ffff8583ffffdad800007a7d;
    assign coff[23  ] = 256'hffff8583ffffdad800007a7d00002528ffff8583ffffdad800007a7d00002528;
    assign coff[24  ] = 256'h00007a7dffffdad8ffff85830000252800007a7dffffdad8ffff858300002528;
    assign coff[25  ] = 256'hffffdad8ffff85830000252800007a7dffffdad8ffff85830000252800007a7d;
    assign coff[26  ] = 256'h00003c57ffff8f1dffffc3a9000070e300003c57ffff8f1dffffc3a9000070e3;
    assign coff[27  ] = 256'hffff8f1dffffc3a9000070e300003c57ffff8f1dffffc3a9000070e300003c57;
    assign coff[28  ] = 256'h000062f2ffffaeccffff9d0e00005134000062f2ffffaeccffff9d0e00005134;
    assign coff[29  ] = 256'hffffaeccffff9d0e00005134000062f2ffffaeccffff9d0e00005134000062f2;
    assign coff[30  ] = 256'h00000c8cffff809efffff37400007f6200000c8cffff809efffff37400007f62;
    assign coff[31  ] = 256'hffff809efffff37400007f6200000c8cffff809efffff37400007f6200000c8c;
    assign coff[32  ] = 256'h00007fd9fffff9b8ffff80270000064800007fd9fffff9b8ffff802700000648;
    assign coff[33  ] = 256'hfffff9b8ffff80270000064800007fd9fffff9b8ffff80270000064800007fd9;
    assign coff[34  ] = 256'h000055f6ffffa129ffffaa0a00005ed7000055f6ffffa129ffffaa0a00005ed7;
    assign coff[35  ] = 256'hffffa129ffffaa0a00005ed7000055f6ffffa129ffffaa0a00005ed7000055f6;
    assign coff[36  ] = 256'h000073b6ffffc946ffff8c4a000036ba000073b6ffffc946ffff8c4a000036ba;
    assign coff[37  ] = 256'hffffc946ffff8c4a000036ba000073b6ffffc946ffff8c4a000036ba000073b6;
    assign coff[38  ] = 256'h00002b1fffff877bffffd4e10000788500002b1fffff877bffffd4e100007885;
    assign coff[39  ] = 256'hffff877bffffd4e10000788500002b1fffff877bffffd4e10000788500002b1f;
    assign coff[40  ] = 256'h00007c2affffe0e6ffff83d600001f1a00007c2affffe0e6ffff83d600001f1a;
    assign coff[41  ] = 256'hffffe0e6ffff83d600001f1a00007c2affffe0e6ffff83d600001f1a00007c2a;
    assign coff[42  ] = 256'h000041ceffff9236ffffbe3200006dca000041ceffff9236ffffbe3200006dca;
    assign coff[43  ] = 256'hffff9236ffffbe3200006dca000041ceffff9236ffffbe3200006dca000041ce;
    assign coff[44  ] = 256'h000066d0ffffb3c0ffff993000004c40000066d0ffffb3c0ffff993000004c40;
    assign coff[45  ] = 256'hffffb3c0ffff993000004c40000066d0ffffb3c0ffff993000004c40000066d0;
    assign coff[46  ] = 256'h000012c8ffff8163ffffed3800007e9d000012c8ffff8163ffffed3800007e9d;
    assign coff[47  ] = 256'hffff8163ffffed3800007e9d000012c8ffff8163ffffed3800007e9d000012c8;
    assign coff[48  ] = 256'h00007e9dffffed38ffff8163000012c800007e9dffffed38ffff8163000012c8;
    assign coff[49  ] = 256'hffffed38ffff8163000012c800007e9dffffed38ffff8163000012c800007e9d;
    assign coff[50  ] = 256'h00004c40ffff9930ffffb3c0000066d000004c40ffff9930ffffb3c0000066d0;
    assign coff[51  ] = 256'hffff9930ffffb3c0000066d000004c40ffff9930ffffb3c0000066d000004c40;
    assign coff[52  ] = 256'h00006dcaffffbe32ffff9236000041ce00006dcaffffbe32ffff9236000041ce;
    assign coff[53  ] = 256'hffffbe32ffff9236000041ce00006dcaffffbe32ffff9236000041ce00006dca;
    assign coff[54  ] = 256'h00001f1affff83d6ffffe0e600007c2a00001f1affff83d6ffffe0e600007c2a;
    assign coff[55  ] = 256'hffff83d6ffffe0e600007c2a00001f1affff83d6ffffe0e600007c2a00001f1a;
    assign coff[56  ] = 256'h00007885ffffd4e1ffff877b00002b1f00007885ffffd4e1ffff877b00002b1f;
    assign coff[57  ] = 256'hffffd4e1ffff877b00002b1f00007885ffffd4e1ffff877b00002b1f00007885;
    assign coff[58  ] = 256'h000036baffff8c4affffc946000073b6000036baffff8c4affffc946000073b6;
    assign coff[59  ] = 256'hffff8c4affffc946000073b6000036baffff8c4affffc946000073b6000036ba;
    assign coff[60  ] = 256'h00005ed7ffffaa0affffa129000055f600005ed7ffffaa0affffa129000055f6;
    assign coff[61  ] = 256'hffffaa0affffa129000055f600005ed7ffffaa0affffa129000055f600005ed7;
    assign coff[62  ] = 256'h00000648ffff8027fffff9b800007fd900000648ffff8027fffff9b800007fd9;
    assign coff[63  ] = 256'hffff8027fffff9b800007fd900000648ffff8027fffff9b800007fd900000648;
    assign coff[64  ] = 256'h00007ff6fffffcdcffff800a0000032400007ff6fffffcdcffff800a00000324;
    assign coff[65  ] = 256'hfffffcdcffff800a0000032400007ff6fffffcdcffff800a0000032400007ff6;
    assign coff[66  ] = 256'h00005843ffffa34cffffa7bd00005cb400005843ffffa34cffffa7bd00005cb4;
    assign coff[67  ] = 256'hffffa34cffffa7bd00005cb400005843ffffa34cffffa7bd00005cb400005843;
    assign coff[68  ] = 256'h00007505ffffcc21ffff8afb000033df00007505ffffcc21ffff8afb000033df;
    assign coff[69  ] = 256'hffffcc21ffff8afb000033df00007505ffffcc21ffff8afb000033df00007505;
    assign coff[70  ] = 256'h00002e11ffff8894ffffd1ef0000776c00002e11ffff8894ffffd1ef0000776c;
    assign coff[71  ] = 256'hffff8894ffffd1ef0000776c00002e11ffff8894ffffd1ef0000776c00002e11;
    assign coff[72  ] = 256'h00007ce4ffffe3f4ffff831c00001c0c00007ce4ffffe3f4ffff831c00001c0c;
    assign coff[73  ] = 256'hffffe3f4ffff831c00001c0c00007ce4ffffe3f4ffff831c00001c0c00007ce4;
    assign coff[74  ] = 256'h0000447bffff93dcffffbb8500006c240000447bffff93dcffffbb8500006c24;
    assign coff[75  ] = 256'hffff93dcffffbb8500006c240000447bffff93dcffffbb8500006c240000447b;
    assign coff[76  ] = 256'h000068a7ffffb64cffff9759000049b4000068a7ffffb64cffff9759000049b4;
    assign coff[77  ] = 256'hffffb64cffff9759000049b4000068a7ffffb64cffff9759000049b4000068a7;
    assign coff[78  ] = 256'h000015e2ffff81e2ffffea1e00007e1e000015e2ffff81e2ffffea1e00007e1e;
    assign coff[79  ] = 256'hffff81e2ffffea1e00007e1e000015e2ffff81e2ffffea1e00007e1e000015e2;
    assign coff[80  ] = 256'h00007f0afffff055ffff80f600000fab00007f0afffff055ffff80f600000fab;
    assign coff[81  ] = 256'hfffff055ffff80f600000fab00007f0afffff055ffff80f600000fab00007f0a;
    assign coff[82  ] = 256'h00004ec0ffff9b17ffffb140000064e900004ec0ffff9b17ffffb140000064e9;
    assign coff[83  ] = 256'hffff9b17ffffb140000064e900004ec0ffff9b17ffffb140000064e900004ec0;
    assign coff[84  ] = 256'h00006f5fffffc0e9ffff90a100003f1700006f5fffffc0e9ffff90a100003f17;
    assign coff[85  ] = 256'hffffc0e9ffff90a100003f1700006f5fffffc0e9ffff90a100003f1700006f5f;
    assign coff[86  ] = 256'h00002224ffff84a3ffffdddc00007b5d00002224ffff84a3ffffdddc00007b5d;
    assign coff[87  ] = 256'hffff84a3ffffdddc00007b5d00002224ffff84a3ffffdddc00007b5d00002224;
    assign coff[88  ] = 256'h0000798affffd7d9ffff8676000028270000798affffd7d9ffff867600002827;
    assign coff[89  ] = 256'hffffd7d9ffff8676000028270000798affffd7d9ffff8676000028270000798a;
    assign coff[90  ] = 256'h0000398dffff8dabffffc673000072550000398dffff8dabffffc67300007255;
    assign coff[91  ] = 256'hffff8dabffffc673000072550000398dffff8dabffffc673000072550000398d;
    assign coff[92  ] = 256'h000060ecffffac65ffff9f140000539b000060ecffffac65ffff9f140000539b;
    assign coff[93  ] = 256'hffffac65ffff9f140000539b000060ecffffac65ffff9f140000539b000060ec;
    assign coff[94  ] = 256'h0000096bffff8059fffff69500007fa70000096bffff8059fffff69500007fa7;
    assign coff[95  ] = 256'hffff8059fffff69500007fa70000096bffff8059fffff69500007fa70000096b;
    assign coff[96  ] = 256'h00007fa7fffff695ffff80590000096b00007fa7fffff695ffff80590000096b;
    assign coff[97  ] = 256'hfffff695ffff80590000096b00007fa7fffff695ffff80590000096b00007fa7;
    assign coff[98  ] = 256'h0000539bffff9f14ffffac65000060ec0000539bffff9f14ffffac65000060ec;
    assign coff[99  ] = 256'hffff9f14ffffac65000060ec0000539bffff9f14ffffac65000060ec0000539b;
    assign coff[100 ] = 256'h00007255ffffc673ffff8dab0000398d00007255ffffc673ffff8dab0000398d;
    assign coff[101 ] = 256'hffffc673ffff8dab0000398d00007255ffffc673ffff8dab0000398d00007255;
    assign coff[102 ] = 256'h00002827ffff8676ffffd7d90000798a00002827ffff8676ffffd7d90000798a;
    assign coff[103 ] = 256'hffff8676ffffd7d90000798a00002827ffff8676ffffd7d90000798a00002827;
    assign coff[104 ] = 256'h00007b5dffffdddcffff84a30000222400007b5dffffdddcffff84a300002224;
    assign coff[105 ] = 256'hffffdddcffff84a30000222400007b5dffffdddcffff84a30000222400007b5d;
    assign coff[106 ] = 256'h00003f17ffff90a1ffffc0e900006f5f00003f17ffff90a1ffffc0e900006f5f;
    assign coff[107 ] = 256'hffff90a1ffffc0e900006f5f00003f17ffff90a1ffffc0e900006f5f00003f17;
    assign coff[108 ] = 256'h000064e9ffffb140ffff9b1700004ec0000064e9ffffb140ffff9b1700004ec0;
    assign coff[109 ] = 256'hffffb140ffff9b1700004ec0000064e9ffffb140ffff9b1700004ec0000064e9;
    assign coff[110 ] = 256'h00000fabffff80f6fffff05500007f0a00000fabffff80f6fffff05500007f0a;
    assign coff[111 ] = 256'hffff80f6fffff05500007f0a00000fabffff80f6fffff05500007f0a00000fab;
    assign coff[112 ] = 256'h00007e1effffea1effff81e2000015e200007e1effffea1effff81e2000015e2;
    assign coff[113 ] = 256'hffffea1effff81e2000015e200007e1effffea1effff81e2000015e200007e1e;
    assign coff[114 ] = 256'h000049b4ffff9759ffffb64c000068a7000049b4ffff9759ffffb64c000068a7;
    assign coff[115 ] = 256'hffff9759ffffb64c000068a7000049b4ffff9759ffffb64c000068a7000049b4;
    assign coff[116 ] = 256'h00006c24ffffbb85ffff93dc0000447b00006c24ffffbb85ffff93dc0000447b;
    assign coff[117 ] = 256'hffffbb85ffff93dc0000447b00006c24ffffbb85ffff93dc0000447b00006c24;
    assign coff[118 ] = 256'h00001c0cffff831cffffe3f400007ce400001c0cffff831cffffe3f400007ce4;
    assign coff[119 ] = 256'hffff831cffffe3f400007ce400001c0cffff831cffffe3f400007ce400001c0c;
    assign coff[120 ] = 256'h0000776cffffd1efffff889400002e110000776cffffd1efffff889400002e11;
    assign coff[121 ] = 256'hffffd1efffff889400002e110000776cffffd1efffff889400002e110000776c;
    assign coff[122 ] = 256'h000033dfffff8afbffffcc2100007505000033dfffff8afbffffcc2100007505;
    assign coff[123 ] = 256'hffff8afbffffcc2100007505000033dfffff8afbffffcc2100007505000033df;
    assign coff[124 ] = 256'h00005cb4ffffa7bdffffa34c0000584300005cb4ffffa7bdffffa34c00005843;
    assign coff[125 ] = 256'hffffa7bdffffa34c0000584300005cb4ffffa7bdffffa34c0000584300005cb4;
    assign coff[126 ] = 256'h00000324ffff800afffffcdc00007ff600000324ffff800afffffcdc00007ff6;
    assign coff[127 ] = 256'hffff800afffffcdc00007ff600000324ffff800afffffcdc00007ff600000324;
    assign coff[128 ] = 256'h00007ffefffffe6effff80020000019200007ffefffffe6effff800200000192;
    assign coff[129 ] = 256'hfffffe6effff80020000019200007ffefffffe6effff80020000019200007ffe;
    assign coff[130 ] = 256'h00005964ffffa463ffffa69c00005b9d00005964ffffa463ffffa69c00005b9d;
    assign coff[131 ] = 256'hffffa463ffffa69c00005b9d00005964ffffa463ffffa69c00005b9d00005964;
    assign coff[132 ] = 256'h000075a6ffffcd92ffff8a5a0000326e000075a6ffffcd92ffff8a5a0000326e;
    assign coff[133 ] = 256'hffffcd92ffff8a5a0000326e000075a6ffffcd92ffff8a5a0000326e000075a6;
    assign coff[134 ] = 256'h00002f87ffff8927ffffd079000076d900002f87ffff8927ffffd079000076d9;
    assign coff[135 ] = 256'hffff8927ffffd079000076d900002f87ffff8927ffffd079000076d900002f87;
    assign coff[136 ] = 256'h00007d3affffe57dffff82c600001a8300007d3affffe57dffff82c600001a83;
    assign coff[137 ] = 256'hffffe57dffff82c600001a8300007d3affffe57dffff82c600001a8300007d3a;
    assign coff[138 ] = 256'h000045cdffff94b5ffffba3300006b4b000045cdffff94b5ffffba3300006b4b;
    assign coff[139 ] = 256'hffff94b5ffffba3300006b4b000045cdffff94b5ffffba3300006b4b000045cd;
    assign coff[140 ] = 256'h0000698cffffb796ffff96740000486a0000698cffffb796ffff96740000486a;
    assign coff[141 ] = 256'hffffb796ffff96740000486a0000698cffffb796ffff96740000486a0000698c;
    assign coff[142 ] = 256'h0000176effff822affffe89200007dd60000176effff822affffe89200007dd6;
    assign coff[143 ] = 256'hffff822affffe89200007dd60000176effff822affffe89200007dd60000176e;
    assign coff[144 ] = 256'h00007f38fffff1e4ffff80c800000e1c00007f38fffff1e4ffff80c800000e1c;
    assign coff[145 ] = 256'hfffff1e4ffff80c800000e1c00007f38fffff1e4ffff80c800000e1c00007f38;
    assign coff[146 ] = 256'h00004ffbffff9c11ffffb005000063ef00004ffbffff9c11ffffb005000063ef;
    assign coff[147 ] = 256'hffff9c11ffffb005000063ef00004ffbffff9c11ffffb005000063ef00004ffb;
    assign coff[148 ] = 256'h00007023ffffc248ffff8fdd00003db800007023ffffc248ffff8fdd00003db8;
    assign coff[149 ] = 256'hffffc248ffff8fdd00003db800007023ffffc248ffff8fdd00003db800007023;
    assign coff[150 ] = 256'h000023a7ffff8511ffffdc5900007aef000023a7ffff8511ffffdc5900007aef;
    assign coff[151 ] = 256'hffff8511ffffdc5900007aef000023a7ffff8511ffffdc5900007aef000023a7;
    assign coff[152 ] = 256'h00007a06ffffd958ffff85fa000026a800007a06ffffd958ffff85fa000026a8;
    assign coff[153 ] = 256'hffffd958ffff85fa000026a800007a06ffffd958ffff85fa000026a800007a06;
    assign coff[154 ] = 256'h00003af3ffff8e62ffffc50d0000719e00003af3ffff8e62ffffc50d0000719e;
    assign coff[155 ] = 256'hffff8e62ffffc50d0000719e00003af3ffff8e62ffffc50d0000719e00003af3;
    assign coff[156 ] = 256'h000061f1ffffad97ffff9e0f00005269000061f1ffffad97ffff9e0f00005269;
    assign coff[157 ] = 256'hffffad97ffff9e0f00005269000061f1ffffad97ffff9e0f00005269000061f1;
    assign coff[158 ] = 256'h00000afbffff8079fffff50500007f8700000afbffff8079fffff50500007f87;
    assign coff[159 ] = 256'hffff8079fffff50500007f8700000afbffff8079fffff50500007f8700000afb;
    assign coff[160 ] = 256'h00007fc2fffff827ffff803e000007d900007fc2fffff827ffff803e000007d9;
    assign coff[161 ] = 256'hfffff827ffff803e000007d900007fc2fffff827ffff803e000007d900007fc2;
    assign coff[162 ] = 256'h000054caffffa01cffffab3600005fe4000054caffffa01cffffab3600005fe4;
    assign coff[163 ] = 256'hffffa01cffffab3600005fe4000054caffffa01cffffab3600005fe4000054ca;
    assign coff[164 ] = 256'h00007308ffffc7dbffff8cf80000382500007308ffffc7dbffff8cf800003825;
    assign coff[165 ] = 256'hffffc7dbffff8cf80000382500007308ffffc7dbffff8cf80000382500007308;
    assign coff[166 ] = 256'h000029a4ffff86f6ffffd65c0000790a000029a4ffff86f6ffffd65c0000790a;
    assign coff[167 ] = 256'hffff86f6ffffd65c0000790a000029a4ffff86f6ffffd65c0000790a000029a4;
    assign coff[168 ] = 256'h00007bc6ffffdf61ffff843a0000209f00007bc6ffffdf61ffff843a0000209f;
    assign coff[169 ] = 256'hffffdf61ffff843a0000209f00007bc6ffffdf61ffff843a0000209f00007bc6;
    assign coff[170 ] = 256'h00004074ffff9169ffffbf8c00006e9700004074ffff9169ffffbf8c00006e97;
    assign coff[171 ] = 256'hffff9169ffffbf8c00006e9700004074ffff9169ffffbf8c00006e9700004074;
    assign coff[172 ] = 256'h000065deffffb27fffff9a2200004d81000065deffffb27fffff9a2200004d81;
    assign coff[173 ] = 256'hffffb27fffff9a2200004d81000065deffffb27fffff9a2200004d81000065de;
    assign coff[174 ] = 256'h0000113affff812affffeec600007ed60000113affff812affffeec600007ed6;
    assign coff[175 ] = 256'hffff812affffeec600007ed60000113affff812affffeec600007ed60000113a;
    assign coff[176 ] = 256'h00007e60ffffebabffff81a00000145500007e60ffffebabffff81a000001455;
    assign coff[177 ] = 256'hffffebabffff81a00000145500007e60ffffebabffff81a00000145500007e60;
    assign coff[178 ] = 256'h00004afbffff9843ffffb505000067bd00004afbffff9843ffffb505000067bd;
    assign coff[179 ] = 256'hffff9843ffffb505000067bd00004afbffff9843ffffb505000067bd00004afb;
    assign coff[180 ] = 256'h00006cf9ffffbcdaffff93070000432600006cf9ffffbcdaffff930700004326;
    assign coff[181 ] = 256'hffffbcdaffff93070000432600006cf9ffffbcdaffff93070000432600006cf9;
    assign coff[182 ] = 256'h00001d93ffff8377ffffe26d00007c8900001d93ffff8377ffffe26d00007c89;
    assign coff[183 ] = 256'hffff8377ffffe26d00007c8900001d93ffff8377ffffe26d00007c8900001d93;
    assign coff[184 ] = 256'h000077fbffffd367ffff880500002c99000077fbffffd367ffff880500002c99;
    assign coff[185 ] = 256'hffffd367ffff880500002c99000077fbffffd367ffff880500002c99000077fb;
    assign coff[186 ] = 256'h0000354effff8ba0ffffcab2000074600000354effff8ba0ffffcab200007460;
    assign coff[187 ] = 256'hffff8ba0ffffcab2000074600000354effff8ba0ffffcab2000074600000354e;
    assign coff[188 ] = 256'h00005dc8ffffa8e2ffffa2380000571e00005dc8ffffa8e2ffffa2380000571e;
    assign coff[189 ] = 256'hffffa8e2ffffa2380000571e00005dc8ffffa8e2ffffa2380000571e00005dc8;
    assign coff[190 ] = 256'h000004b6ffff8016fffffb4a00007fea000004b6ffff8016fffffb4a00007fea;
    assign coff[191 ] = 256'hffff8016fffffb4a00007fea000004b6ffff8016fffffb4a00007fea000004b6;
    assign coff[192 ] = 256'h00007feafffffb4affff8016000004b600007feafffffb4affff8016000004b6;
    assign coff[193 ] = 256'hfffffb4affff8016000004b600007feafffffb4affff8016000004b600007fea;
    assign coff[194 ] = 256'h0000571effffa238ffffa8e200005dc80000571effffa238ffffa8e200005dc8;
    assign coff[195 ] = 256'hffffa238ffffa8e200005dc80000571effffa238ffffa8e200005dc80000571e;
    assign coff[196 ] = 256'h00007460ffffcab2ffff8ba00000354e00007460ffffcab2ffff8ba00000354e;
    assign coff[197 ] = 256'hffffcab2ffff8ba00000354e00007460ffffcab2ffff8ba00000354e00007460;
    assign coff[198 ] = 256'h00002c99ffff8805ffffd367000077fb00002c99ffff8805ffffd367000077fb;
    assign coff[199 ] = 256'hffff8805ffffd367000077fb00002c99ffff8805ffffd367000077fb00002c99;
    assign coff[200 ] = 256'h00007c89ffffe26dffff837700001d9300007c89ffffe26dffff837700001d93;
    assign coff[201 ] = 256'hffffe26dffff837700001d9300007c89ffffe26dffff837700001d9300007c89;
    assign coff[202 ] = 256'h00004326ffff9307ffffbcda00006cf900004326ffff9307ffffbcda00006cf9;
    assign coff[203 ] = 256'hffff9307ffffbcda00006cf900004326ffff9307ffffbcda00006cf900004326;
    assign coff[204 ] = 256'h000067bdffffb505ffff984300004afb000067bdffffb505ffff984300004afb;
    assign coff[205 ] = 256'hffffb505ffff984300004afb000067bdffffb505ffff984300004afb000067bd;
    assign coff[206 ] = 256'h00001455ffff81a0ffffebab00007e6000001455ffff81a0ffffebab00007e60;
    assign coff[207 ] = 256'hffff81a0ffffebab00007e6000001455ffff81a0ffffebab00007e6000001455;
    assign coff[208 ] = 256'h00007ed6ffffeec6ffff812a0000113a00007ed6ffffeec6ffff812a0000113a;
    assign coff[209 ] = 256'hffffeec6ffff812a0000113a00007ed6ffffeec6ffff812a0000113a00007ed6;
    assign coff[210 ] = 256'h00004d81ffff9a22ffffb27f000065de00004d81ffff9a22ffffb27f000065de;
    assign coff[211 ] = 256'hffff9a22ffffb27f000065de00004d81ffff9a22ffffb27f000065de00004d81;
    assign coff[212 ] = 256'h00006e97ffffbf8cffff91690000407400006e97ffffbf8cffff916900004074;
    assign coff[213 ] = 256'hffffbf8cffff91690000407400006e97ffffbf8cffff91690000407400006e97;
    assign coff[214 ] = 256'h0000209fffff843affffdf6100007bc60000209fffff843affffdf6100007bc6;
    assign coff[215 ] = 256'hffff843affffdf6100007bc60000209fffff843affffdf6100007bc60000209f;
    assign coff[216 ] = 256'h0000790affffd65cffff86f6000029a40000790affffd65cffff86f6000029a4;
    assign coff[217 ] = 256'hffffd65cffff86f6000029a40000790affffd65cffff86f6000029a40000790a;
    assign coff[218 ] = 256'h00003825ffff8cf8ffffc7db0000730800003825ffff8cf8ffffc7db00007308;
    assign coff[219 ] = 256'hffff8cf8ffffc7db0000730800003825ffff8cf8ffffc7db0000730800003825;
    assign coff[220 ] = 256'h00005fe4ffffab36ffffa01c000054ca00005fe4ffffab36ffffa01c000054ca;
    assign coff[221 ] = 256'hffffab36ffffa01c000054ca00005fe4ffffab36ffffa01c000054ca00005fe4;
    assign coff[222 ] = 256'h000007d9ffff803efffff82700007fc2000007d9ffff803efffff82700007fc2;
    assign coff[223 ] = 256'hffff803efffff82700007fc2000007d9ffff803efffff82700007fc2000007d9;
    assign coff[224 ] = 256'h00007f87fffff505ffff807900000afb00007f87fffff505ffff807900000afb;
    assign coff[225 ] = 256'hfffff505ffff807900000afb00007f87fffff505ffff807900000afb00007f87;
    assign coff[226 ] = 256'h00005269ffff9e0fffffad97000061f100005269ffff9e0fffffad97000061f1;
    assign coff[227 ] = 256'hffff9e0fffffad97000061f100005269ffff9e0fffffad97000061f100005269;
    assign coff[228 ] = 256'h0000719effffc50dffff8e6200003af30000719effffc50dffff8e6200003af3;
    assign coff[229 ] = 256'hffffc50dffff8e6200003af30000719effffc50dffff8e6200003af30000719e;
    assign coff[230 ] = 256'h000026a8ffff85faffffd95800007a06000026a8ffff85faffffd95800007a06;
    assign coff[231 ] = 256'hffff85faffffd95800007a06000026a8ffff85faffffd95800007a06000026a8;
    assign coff[232 ] = 256'h00007aefffffdc59ffff8511000023a700007aefffffdc59ffff8511000023a7;
    assign coff[233 ] = 256'hffffdc59ffff8511000023a700007aefffffdc59ffff8511000023a700007aef;
    assign coff[234 ] = 256'h00003db8ffff8fddffffc2480000702300003db8ffff8fddffffc24800007023;
    assign coff[235 ] = 256'hffff8fddffffc2480000702300003db8ffff8fddffffc2480000702300003db8;
    assign coff[236 ] = 256'h000063efffffb005ffff9c1100004ffb000063efffffb005ffff9c1100004ffb;
    assign coff[237 ] = 256'hffffb005ffff9c1100004ffb000063efffffb005ffff9c1100004ffb000063ef;
    assign coff[238 ] = 256'h00000e1cffff80c8fffff1e400007f3800000e1cffff80c8fffff1e400007f38;
    assign coff[239 ] = 256'hffff80c8fffff1e400007f3800000e1cffff80c8fffff1e400007f3800000e1c;
    assign coff[240 ] = 256'h00007dd6ffffe892ffff822a0000176e00007dd6ffffe892ffff822a0000176e;
    assign coff[241 ] = 256'hffffe892ffff822a0000176e00007dd6ffffe892ffff822a0000176e00007dd6;
    assign coff[242 ] = 256'h0000486affff9674ffffb7960000698c0000486affff9674ffffb7960000698c;
    assign coff[243 ] = 256'hffff9674ffffb7960000698c0000486affff9674ffffb7960000698c0000486a;
    assign coff[244 ] = 256'h00006b4bffffba33ffff94b5000045cd00006b4bffffba33ffff94b5000045cd;
    assign coff[245 ] = 256'hffffba33ffff94b5000045cd00006b4bffffba33ffff94b5000045cd00006b4b;
    assign coff[246 ] = 256'h00001a83ffff82c6ffffe57d00007d3a00001a83ffff82c6ffffe57d00007d3a;
    assign coff[247 ] = 256'hffff82c6ffffe57d00007d3a00001a83ffff82c6ffffe57d00007d3a00001a83;
    assign coff[248 ] = 256'h000076d9ffffd079ffff892700002f87000076d9ffffd079ffff892700002f87;
    assign coff[249 ] = 256'hffffd079ffff892700002f87000076d9ffffd079ffff892700002f87000076d9;
    assign coff[250 ] = 256'h0000326effff8a5affffcd92000075a60000326effff8a5affffcd92000075a6;
    assign coff[251 ] = 256'hffff8a5affffcd92000075a60000326effff8a5affffcd92000075a60000326e;
    assign coff[252 ] = 256'h00005b9dffffa69cffffa4630000596400005b9dffffa69cffffa46300005964;
    assign coff[253 ] = 256'hffffa69cffffa4630000596400005b9dffffa69cffffa4630000596400005b9d;
    assign coff[254 ] = 256'h00000192ffff8002fffffe6e00007ffe00000192ffff8002fffffe6e00007ffe;
    assign coff[255 ] = 256'hffff8002fffffe6e00007ffe00000192ffff8002fffffe6e00007ffe00000192;
    assign coff[256 ] = 256'h00007fffffffff37ffff8001000000c900007fffffffff37ffff8001000000c9;
    assign coff[257 ] = 256'hffffff37ffff8001000000c900007fffffffff37ffff8001000000c900007fff;
    assign coff[258 ] = 256'h000059f4ffffa4f0ffffa60c00005b10000059f4ffffa4f0ffffa60c00005b10;
    assign coff[259 ] = 256'hffffa4f0ffffa60c00005b10000059f4ffffa4f0ffffa60c00005b10000059f4;
    assign coff[260 ] = 256'h000075f4ffffce4bffff8a0c000031b5000075f4ffffce4bffff8a0c000031b5;
    assign coff[261 ] = 256'hffffce4bffff8a0c000031b5000075f4ffffce4bffff8a0c000031b5000075f4;
    assign coff[262 ] = 256'h00003042ffff8972ffffcfbe0000768e00003042ffff8972ffffcfbe0000768e;
    assign coff[263 ] = 256'hffff8972ffffcfbe0000768e00003042ffff8972ffffcfbe0000768e00003042;
    assign coff[264 ] = 256'h00007d63ffffe642ffff829d000019be00007d63ffffe642ffff829d000019be;
    assign coff[265 ] = 256'hffffe642ffff829d000019be00007d63ffffe642ffff829d000019be00007d63;
    assign coff[266 ] = 256'h00004675ffff9523ffffb98b00006add00004675ffff9523ffffb98b00006add;
    assign coff[267 ] = 256'hffff9523ffffb98b00006add00004675ffff9523ffffb98b00006add00004675;
    assign coff[268 ] = 256'h000069fdffffb83cffff9603000047c4000069fdffffb83cffff9603000047c4;
    assign coff[269 ] = 256'hffffb83cffff9603000047c4000069fdffffb83cffff9603000047c4000069fd;
    assign coff[270 ] = 256'h00001833ffff824fffffe7cd00007db100001833ffff824fffffe7cd00007db1;
    assign coff[271 ] = 256'hffff824fffffe7cd00007db100001833ffff824fffffe7cd00007db100001833;
    assign coff[272 ] = 256'h00007f4efffff2acffff80b200000d5400007f4efffff2acffff80b200000d54;
    assign coff[273 ] = 256'hfffff2acffff80b200000d5400007f4efffff2acffff80b200000d5400007f4e;
    assign coff[274 ] = 256'h00005098ffff9c8fffffaf680000637100005098ffff9c8fffffaf6800006371;
    assign coff[275 ] = 256'hffff9c8fffffaf680000637100005098ffff9c8fffffaf680000637100005098;
    assign coff[276 ] = 256'h00007083ffffc2f8ffff8f7d00003d0800007083ffffc2f8ffff8f7d00003d08;
    assign coff[277 ] = 256'hffffc2f8ffff8f7d00003d0800007083ffffc2f8ffff8f7d00003d0800007083;
    assign coff[278 ] = 256'h00002467ffff8549ffffdb9900007ab700002467ffff8549ffffdb9900007ab7;
    assign coff[279 ] = 256'hffff8549ffffdb9900007ab700002467ffff8549ffffdb9900007ab700002467;
    assign coff[280 ] = 256'h00007a42ffffda18ffff85be000025e800007a42ffffda18ffff85be000025e8;
    assign coff[281 ] = 256'hffffda18ffff85be000025e800007a42ffffda18ffff85be000025e800007a42;
    assign coff[282 ] = 256'h00003ba5ffff8ebfffffc45b0000714100003ba5ffff8ebfffffc45b00007141;
    assign coff[283 ] = 256'hffff8ebfffffc45b0000714100003ba5ffff8ebfffffc45b0000714100003ba5;
    assign coff[284 ] = 256'h00006272ffffae31ffff9d8e000051cf00006272ffffae31ffff9d8e000051cf;
    assign coff[285 ] = 256'hffffae31ffff9d8e000051cf00006272ffffae31ffff9d8e000051cf00006272;
    assign coff[286 ] = 256'h00000bc4ffff808bfffff43c00007f7500000bc4ffff808bfffff43c00007f75;
    assign coff[287 ] = 256'hffff808bfffff43c00007f7500000bc4ffff808bfffff43c00007f7500000bc4;
    assign coff[288 ] = 256'h00007fcefffff8efffff80320000071100007fcefffff8efffff803200000711;
    assign coff[289 ] = 256'hfffff8efffff80320000071100007fcefffff8efffff80320000071100007fce;
    assign coff[290 ] = 256'h00005560ffffa0a2ffffaaa000005f5e00005560ffffa0a2ffffaaa000005f5e;
    assign coff[291 ] = 256'hffffa0a2ffffaaa000005f5e00005560ffffa0a2ffffaaa000005f5e00005560;
    assign coff[292 ] = 256'h0000735fffffc890ffff8ca1000037700000735fffffc890ffff8ca100003770;
    assign coff[293 ] = 256'hffffc890ffff8ca1000037700000735fffffc890ffff8ca1000037700000735f;
    assign coff[294 ] = 256'h00002a62ffff8738ffffd59e000078c800002a62ffff8738ffffd59e000078c8;
    assign coff[295 ] = 256'hffff8738ffffd59e000078c800002a62ffff8738ffffd59e000078c800002a62;
    assign coff[296 ] = 256'h00007bf9ffffe023ffff840700001fdd00007bf9ffffe023ffff840700001fdd;
    assign coff[297 ] = 256'hffffe023ffff840700001fdd00007bf9ffffe023ffff840700001fdd00007bf9;
    assign coff[298 ] = 256'h00004121ffff91cfffffbedf00006e3100004121ffff91cfffffbedf00006e31;
    assign coff[299 ] = 256'hffff91cfffffbedf00006e3100004121ffff91cfffffbedf00006e3100004121;
    assign coff[300 ] = 256'h00006657ffffb31fffff99a900004ce100006657ffffb31fffff99a900004ce1;
    assign coff[301 ] = 256'hffffb31fffff99a900004ce100006657ffffb31fffff99a900004ce100006657;
    assign coff[302 ] = 256'h00001201ffff8146ffffedff00007eba00001201ffff8146ffffedff00007eba;
    assign coff[303 ] = 256'hffff8146ffffedff00007eba00001201ffff8146ffffedff00007eba00001201;
    assign coff[304 ] = 256'h00007e7fffffec71ffff81810000138f00007e7fffffec71ffff81810000138f;
    assign coff[305 ] = 256'hffffec71ffff81810000138f00007e7fffffec71ffff81810000138f00007e7f;
    assign coff[306 ] = 256'h00004b9effff98b9ffffb4620000674700004b9effff98b9ffffb46200006747;
    assign coff[307 ] = 256'hffff98b9ffffb4620000674700004b9effff98b9ffffb4620000674700004b9e;
    assign coff[308 ] = 256'h00006d62ffffbd86ffff929e0000427a00006d62ffffbd86ffff929e0000427a;
    assign coff[309 ] = 256'hffffbd86ffff929e0000427a00006d62ffffbd86ffff929e0000427a00006d62;
    assign coff[310 ] = 256'h00001e57ffff83a6ffffe1a900007c5a00001e57ffff83a6ffffe1a900007c5a;
    assign coff[311 ] = 256'hffff83a6ffffe1a900007c5a00001e57ffff83a6ffffe1a900007c5a00001e57;
    assign coff[312 ] = 256'h00007840ffffd424ffff87c000002bdc00007840ffffd424ffff87c000002bdc;
    assign coff[313 ] = 256'hffffd424ffff87c000002bdc00007840ffffd424ffff87c000002bdc00007840;
    assign coff[314 ] = 256'h00003604ffff8bf5ffffc9fc0000740b00003604ffff8bf5ffffc9fc0000740b;
    assign coff[315 ] = 256'hffff8bf5ffffc9fc0000740b00003604ffff8bf5ffffc9fc0000740b00003604;
    assign coff[316 ] = 256'h00005e50ffffa976ffffa1b00000568a00005e50ffffa976ffffa1b00000568a;
    assign coff[317 ] = 256'hffffa976ffffa1b00000568a00005e50ffffa976ffffa1b00000568a00005e50;
    assign coff[318 ] = 256'h0000057fffff801efffffa8100007fe20000057fffff801efffffa8100007fe2;
    assign coff[319 ] = 256'hffff801efffffa8100007fe20000057fffff801efffffa8100007fe20000057f;
    assign coff[320 ] = 256'h00007ff1fffffc13ffff800f000003ed00007ff1fffffc13ffff800f000003ed;
    assign coff[321 ] = 256'hfffffc13ffff800f000003ed00007ff1fffffc13ffff800f000003ed00007ff1;
    assign coff[322 ] = 256'h000057b1ffffa2c2ffffa84f00005d3e000057b1ffffa2c2ffffa84f00005d3e;
    assign coff[323 ] = 256'hffffa2c2ffffa84f00005d3e000057b1ffffa2c2ffffa84f00005d3e000057b1;
    assign coff[324 ] = 256'h000074b3ffffcb69ffff8b4d00003497000074b3ffffcb69ffff8b4d00003497;
    assign coff[325 ] = 256'hffffcb69ffff8b4d00003497000074b3ffffcb69ffff8b4d00003497000074b3;
    assign coff[326 ] = 256'h00002d55ffff884cffffd2ab000077b400002d55ffff884cffffd2ab000077b4;
    assign coff[327 ] = 256'hffff884cffffd2ab000077b400002d55ffff884cffffd2ab000077b400002d55;
    assign coff[328 ] = 256'h00007cb7ffffe330ffff834900001cd000007cb7ffffe330ffff834900001cd0;
    assign coff[329 ] = 256'hffffe330ffff834900001cd000007cb7ffffe330ffff834900001cd000007cb7;
    assign coff[330 ] = 256'h000043d1ffff9371ffffbc2f00006c8f000043d1ffff9371ffffbc2f00006c8f;
    assign coff[331 ] = 256'hffff9371ffffbc2f00006c8f000043d1ffff9371ffffbc2f00006c8f000043d1;
    assign coff[332 ] = 256'h00006832ffffb5a8ffff97ce00004a5800006832ffffb5a8ffff97ce00004a58;
    assign coff[333 ] = 256'hffffb5a8ffff97ce00004a5800006832ffffb5a8ffff97ce00004a5800006832;
    assign coff[334 ] = 256'h0000151cffff81c1ffffeae400007e3f0000151cffff81c1ffffeae400007e3f;
    assign coff[335 ] = 256'hffff81c1ffffeae400007e3f0000151cffff81c1ffffeae400007e3f0000151c;
    assign coff[336 ] = 256'h00007ef0ffffef8dffff81100000107300007ef0ffffef8dffff811000001073;
    assign coff[337 ] = 256'hffffef8dffff81100000107300007ef0ffffef8dffff81100000107300007ef0;
    assign coff[338 ] = 256'h00004e21ffff9a9cffffb1df0000656400004e21ffff9a9cffffb1df00006564;
    assign coff[339 ] = 256'hffff9a9cffffb1df0000656400004e21ffff9a9cffffb1df0000656400004e21;
    assign coff[340 ] = 256'h00006efbffffc03affff910500003fc600006efbffffc03affff910500003fc6;
    assign coff[341 ] = 256'hffffc03affff910500003fc600006efbffffc03affff910500003fc600006efb;
    assign coff[342 ] = 256'h00002162ffff846effffde9e00007b9200002162ffff846effffde9e00007b92;
    assign coff[343 ] = 256'hffff846effffde9e00007b9200002162ffff846effffde9e00007b9200002162;
    assign coff[344 ] = 256'h0000794affffd71bffff86b6000028e50000794affffd71bffff86b6000028e5;
    assign coff[345 ] = 256'hffffd71bffff86b6000028e50000794affffd71bffff86b6000028e50000794a;
    assign coff[346 ] = 256'h000038d9ffff8d51ffffc727000072af000038d9ffff8d51ffffc727000072af;
    assign coff[347 ] = 256'hffff8d51ffffc727000072af000038d9ffff8d51ffffc727000072af000038d9;
    assign coff[348 ] = 256'h00006068ffffabcdffff9f980000543300006068ffffabcdffff9f9800005433;
    assign coff[349 ] = 256'hffffabcdffff9f980000543300006068ffffabcdffff9f980000543300006068;
    assign coff[350 ] = 256'h000008a2ffff804bfffff75e00007fb5000008a2ffff804bfffff75e00007fb5;
    assign coff[351 ] = 256'hffff804bfffff75e00007fb5000008a2ffff804bfffff75e00007fb5000008a2;
    assign coff[352 ] = 256'h00007f98fffff5cdffff806800000a3300007f98fffff5cdffff806800000a33;
    assign coff[353 ] = 256'hfffff5cdffff806800000a3300007f98fffff5cdffff806800000a3300007f98;
    assign coff[354 ] = 256'h00005303ffff9e91ffffacfd0000616f00005303ffff9e91ffffacfd0000616f;
    assign coff[355 ] = 256'hffff9e91ffffacfd0000616f00005303ffff9e91ffffacfd0000616f00005303;
    assign coff[356 ] = 256'h000071faffffc5c0ffff8e0600003a40000071faffffc5c0ffff8e0600003a40;
    assign coff[357 ] = 256'hffffc5c0ffff8e0600003a40000071faffffc5c0ffff8e0600003a40000071fa;
    assign coff[358 ] = 256'h00002768ffff8637ffffd898000079c900002768ffff8637ffffd898000079c9;
    assign coff[359 ] = 256'hffff8637ffffd898000079c900002768ffff8637ffffd898000079c900002768;
    assign coff[360 ] = 256'h00007b27ffffdd1bffff84d9000022e500007b27ffffdd1bffff84d9000022e5;
    assign coff[361 ] = 256'hffffdd1bffff84d9000022e500007b27ffffdd1bffff84d9000022e500007b27;
    assign coff[362 ] = 256'h00003e68ffff903effffc19800006fc200003e68ffff903effffc19800006fc2;
    assign coff[363 ] = 256'hffff903effffc19800006fc200003e68ffff903effffc19800006fc200003e68;
    assign coff[364 ] = 256'h0000646cffffb0a2ffff9b9400004f5e0000646cffffb0a2ffff9b9400004f5e;
    assign coff[365 ] = 256'hffffb0a2ffff9b9400004f5e0000646cffffb0a2ffff9b9400004f5e0000646c;
    assign coff[366 ] = 256'h00000ee4ffff80defffff11c00007f2200000ee4ffff80defffff11c00007f22;
    assign coff[367 ] = 256'hffff80defffff11c00007f2200000ee4ffff80defffff11c00007f2200000ee4;
    assign coff[368 ] = 256'h00007dfbffffe958ffff8205000016a800007dfbffffe958ffff8205000016a8;
    assign coff[369 ] = 256'hffffe958ffff8205000016a800007dfbffffe958ffff8205000016a800007dfb;
    assign coff[370 ] = 256'h0000490fffff96e6ffffb6f10000691a0000490fffff96e6ffffb6f10000691a;
    assign coff[371 ] = 256'hffff96e6ffffb6f10000691a0000490fffff96e6ffffb6f10000691a0000490f;
    assign coff[372 ] = 256'h00006bb8ffffbadcffff94480000452400006bb8ffffbadcffff944800004524;
    assign coff[373 ] = 256'hffffbadcffff94480000452400006bb8ffffbadcffff94480000452400006bb8;
    assign coff[374 ] = 256'h00001b47ffff82f1ffffe4b900007d0f00001b47ffff82f1ffffe4b900007d0f;
    assign coff[375 ] = 256'hffff82f1ffffe4b900007d0f00001b47ffff82f1ffffe4b900007d0f00001b47;
    assign coff[376 ] = 256'h00007723ffffd134ffff88dd00002ecc00007723ffffd134ffff88dd00002ecc;
    assign coff[377 ] = 256'hffffd134ffff88dd00002ecc00007723ffffd134ffff88dd00002ecc00007723;
    assign coff[378 ] = 256'h00003327ffff8aaaffffccd90000755600003327ffff8aaaffffccd900007556;
    assign coff[379 ] = 256'hffff8aaaffffccd90000755600003327ffff8aaaffffccd90000755600003327;
    assign coff[380 ] = 256'h00005c29ffffa72cffffa3d7000058d400005c29ffffa72cffffa3d7000058d4;
    assign coff[381 ] = 256'hffffa72cffffa3d7000058d400005c29ffffa72cffffa3d7000058d400005c29;
    assign coff[382 ] = 256'h0000025bffff8006fffffda500007ffa0000025bffff8006fffffda500007ffa;
    assign coff[383 ] = 256'hffff8006fffffda500007ffa0000025bffff8006fffffda500007ffa0000025b;
    assign coff[384 ] = 256'h00007ffafffffda5ffff80060000025b00007ffafffffda5ffff80060000025b;
    assign coff[385 ] = 256'hfffffda5ffff80060000025b00007ffafffffda5ffff80060000025b00007ffa;
    assign coff[386 ] = 256'h000058d4ffffa3d7ffffa72c00005c29000058d4ffffa3d7ffffa72c00005c29;
    assign coff[387 ] = 256'hffffa3d7ffffa72c00005c29000058d4ffffa3d7ffffa72c00005c29000058d4;
    assign coff[388 ] = 256'h00007556ffffccd9ffff8aaa0000332700007556ffffccd9ffff8aaa00003327;
    assign coff[389 ] = 256'hffffccd9ffff8aaa0000332700007556ffffccd9ffff8aaa0000332700007556;
    assign coff[390 ] = 256'h00002eccffff88ddffffd1340000772300002eccffff88ddffffd13400007723;
    assign coff[391 ] = 256'hffff88ddffffd1340000772300002eccffff88ddffffd1340000772300002ecc;
    assign coff[392 ] = 256'h00007d0fffffe4b9ffff82f100001b4700007d0fffffe4b9ffff82f100001b47;
    assign coff[393 ] = 256'hffffe4b9ffff82f100001b4700007d0fffffe4b9ffff82f100001b4700007d0f;
    assign coff[394 ] = 256'h00004524ffff9448ffffbadc00006bb800004524ffff9448ffffbadc00006bb8;
    assign coff[395 ] = 256'hffff9448ffffbadc00006bb800004524ffff9448ffffbadc00006bb800004524;
    assign coff[396 ] = 256'h0000691affffb6f1ffff96e60000490f0000691affffb6f1ffff96e60000490f;
    assign coff[397 ] = 256'hffffb6f1ffff96e60000490f0000691affffb6f1ffff96e60000490f0000691a;
    assign coff[398 ] = 256'h000016a8ffff8205ffffe95800007dfb000016a8ffff8205ffffe95800007dfb;
    assign coff[399 ] = 256'hffff8205ffffe95800007dfb000016a8ffff8205ffffe95800007dfb000016a8;
    assign coff[400 ] = 256'h00007f22fffff11cffff80de00000ee400007f22fffff11cffff80de00000ee4;
    assign coff[401 ] = 256'hfffff11cffff80de00000ee400007f22fffff11cffff80de00000ee400007f22;
    assign coff[402 ] = 256'h00004f5effff9b94ffffb0a20000646c00004f5effff9b94ffffb0a20000646c;
    assign coff[403 ] = 256'hffff9b94ffffb0a20000646c00004f5effff9b94ffffb0a20000646c00004f5e;
    assign coff[404 ] = 256'h00006fc2ffffc198ffff903e00003e6800006fc2ffffc198ffff903e00003e68;
    assign coff[405 ] = 256'hffffc198ffff903e00003e6800006fc2ffffc198ffff903e00003e6800006fc2;
    assign coff[406 ] = 256'h000022e5ffff84d9ffffdd1b00007b27000022e5ffff84d9ffffdd1b00007b27;
    assign coff[407 ] = 256'hffff84d9ffffdd1b00007b27000022e5ffff84d9ffffdd1b00007b27000022e5;
    assign coff[408 ] = 256'h000079c9ffffd898ffff863700002768000079c9ffffd898ffff863700002768;
    assign coff[409 ] = 256'hffffd898ffff863700002768000079c9ffffd898ffff863700002768000079c9;
    assign coff[410 ] = 256'h00003a40ffff8e06ffffc5c0000071fa00003a40ffff8e06ffffc5c0000071fa;
    assign coff[411 ] = 256'hffff8e06ffffc5c0000071fa00003a40ffff8e06ffffc5c0000071fa00003a40;
    assign coff[412 ] = 256'h0000616fffffacfdffff9e91000053030000616fffffacfdffff9e9100005303;
    assign coff[413 ] = 256'hffffacfdffff9e91000053030000616fffffacfdffff9e91000053030000616f;
    assign coff[414 ] = 256'h00000a33ffff8068fffff5cd00007f9800000a33ffff8068fffff5cd00007f98;
    assign coff[415 ] = 256'hffff8068fffff5cd00007f9800000a33ffff8068fffff5cd00007f9800000a33;
    assign coff[416 ] = 256'h00007fb5fffff75effff804b000008a200007fb5fffff75effff804b000008a2;
    assign coff[417 ] = 256'hfffff75effff804b000008a200007fb5fffff75effff804b000008a200007fb5;
    assign coff[418 ] = 256'h00005433ffff9f98ffffabcd0000606800005433ffff9f98ffffabcd00006068;
    assign coff[419 ] = 256'hffff9f98ffffabcd0000606800005433ffff9f98ffffabcd0000606800005433;
    assign coff[420 ] = 256'h000072afffffc727ffff8d51000038d9000072afffffc727ffff8d51000038d9;
    assign coff[421 ] = 256'hffffc727ffff8d51000038d9000072afffffc727ffff8d51000038d9000072af;
    assign coff[422 ] = 256'h000028e5ffff86b6ffffd71b0000794a000028e5ffff86b6ffffd71b0000794a;
    assign coff[423 ] = 256'hffff86b6ffffd71b0000794a000028e5ffff86b6ffffd71b0000794a000028e5;
    assign coff[424 ] = 256'h00007b92ffffde9effff846e0000216200007b92ffffde9effff846e00002162;
    assign coff[425 ] = 256'hffffde9effff846e0000216200007b92ffffde9effff846e0000216200007b92;
    assign coff[426 ] = 256'h00003fc6ffff9105ffffc03a00006efb00003fc6ffff9105ffffc03a00006efb;
    assign coff[427 ] = 256'hffff9105ffffc03a00006efb00003fc6ffff9105ffffc03a00006efb00003fc6;
    assign coff[428 ] = 256'h00006564ffffb1dfffff9a9c00004e2100006564ffffb1dfffff9a9c00004e21;
    assign coff[429 ] = 256'hffffb1dfffff9a9c00004e2100006564ffffb1dfffff9a9c00004e2100006564;
    assign coff[430 ] = 256'h00001073ffff8110ffffef8d00007ef000001073ffff8110ffffef8d00007ef0;
    assign coff[431 ] = 256'hffff8110ffffef8d00007ef000001073ffff8110ffffef8d00007ef000001073;
    assign coff[432 ] = 256'h00007e3fffffeae4ffff81c10000151c00007e3fffffeae4ffff81c10000151c;
    assign coff[433 ] = 256'hffffeae4ffff81c10000151c00007e3fffffeae4ffff81c10000151c00007e3f;
    assign coff[434 ] = 256'h00004a58ffff97ceffffb5a80000683200004a58ffff97ceffffb5a800006832;
    assign coff[435 ] = 256'hffff97ceffffb5a80000683200004a58ffff97ceffffb5a80000683200004a58;
    assign coff[436 ] = 256'h00006c8fffffbc2fffff9371000043d100006c8fffffbc2fffff9371000043d1;
    assign coff[437 ] = 256'hffffbc2fffff9371000043d100006c8fffffbc2fffff9371000043d100006c8f;
    assign coff[438 ] = 256'h00001cd0ffff8349ffffe33000007cb700001cd0ffff8349ffffe33000007cb7;
    assign coff[439 ] = 256'hffff8349ffffe33000007cb700001cd0ffff8349ffffe33000007cb700001cd0;
    assign coff[440 ] = 256'h000077b4ffffd2abffff884c00002d55000077b4ffffd2abffff884c00002d55;
    assign coff[441 ] = 256'hffffd2abffff884c00002d55000077b4ffffd2abffff884c00002d55000077b4;
    assign coff[442 ] = 256'h00003497ffff8b4dffffcb69000074b300003497ffff8b4dffffcb69000074b3;
    assign coff[443 ] = 256'hffff8b4dffffcb69000074b300003497ffff8b4dffffcb69000074b300003497;
    assign coff[444 ] = 256'h00005d3effffa84fffffa2c2000057b100005d3effffa84fffffa2c2000057b1;
    assign coff[445 ] = 256'hffffa84fffffa2c2000057b100005d3effffa84fffffa2c2000057b100005d3e;
    assign coff[446 ] = 256'h000003edffff800ffffffc1300007ff1000003edffff800ffffffc1300007ff1;
    assign coff[447 ] = 256'hffff800ffffffc1300007ff1000003edffff800ffffffc1300007ff1000003ed;
    assign coff[448 ] = 256'h00007fe2fffffa81ffff801e0000057f00007fe2fffffa81ffff801e0000057f;
    assign coff[449 ] = 256'hfffffa81ffff801e0000057f00007fe2fffffa81ffff801e0000057f00007fe2;
    assign coff[450 ] = 256'h0000568affffa1b0ffffa97600005e500000568affffa1b0ffffa97600005e50;
    assign coff[451 ] = 256'hffffa1b0ffffa97600005e500000568affffa1b0ffffa97600005e500000568a;
    assign coff[452 ] = 256'h0000740bffffc9fcffff8bf5000036040000740bffffc9fcffff8bf500003604;
    assign coff[453 ] = 256'hffffc9fcffff8bf5000036040000740bffffc9fcffff8bf5000036040000740b;
    assign coff[454 ] = 256'h00002bdcffff87c0ffffd4240000784000002bdcffff87c0ffffd42400007840;
    assign coff[455 ] = 256'hffff87c0ffffd4240000784000002bdcffff87c0ffffd4240000784000002bdc;
    assign coff[456 ] = 256'h00007c5affffe1a9ffff83a600001e5700007c5affffe1a9ffff83a600001e57;
    assign coff[457 ] = 256'hffffe1a9ffff83a600001e5700007c5affffe1a9ffff83a600001e5700007c5a;
    assign coff[458 ] = 256'h0000427affff929effffbd8600006d620000427affff929effffbd8600006d62;
    assign coff[459 ] = 256'hffff929effffbd8600006d620000427affff929effffbd8600006d620000427a;
    assign coff[460 ] = 256'h00006747ffffb462ffff98b900004b9e00006747ffffb462ffff98b900004b9e;
    assign coff[461 ] = 256'hffffb462ffff98b900004b9e00006747ffffb462ffff98b900004b9e00006747;
    assign coff[462 ] = 256'h0000138fffff8181ffffec7100007e7f0000138fffff8181ffffec7100007e7f;
    assign coff[463 ] = 256'hffff8181ffffec7100007e7f0000138fffff8181ffffec7100007e7f0000138f;
    assign coff[464 ] = 256'h00007ebaffffedffffff81460000120100007ebaffffedffffff814600001201;
    assign coff[465 ] = 256'hffffedffffff81460000120100007ebaffffedffffff81460000120100007eba;
    assign coff[466 ] = 256'h00004ce1ffff99a9ffffb31f0000665700004ce1ffff99a9ffffb31f00006657;
    assign coff[467 ] = 256'hffff99a9ffffb31f0000665700004ce1ffff99a9ffffb31f0000665700004ce1;
    assign coff[468 ] = 256'h00006e31ffffbedfffff91cf0000412100006e31ffffbedfffff91cf00004121;
    assign coff[469 ] = 256'hffffbedfffff91cf0000412100006e31ffffbedfffff91cf0000412100006e31;
    assign coff[470 ] = 256'h00001fddffff8407ffffe02300007bf900001fddffff8407ffffe02300007bf9;
    assign coff[471 ] = 256'hffff8407ffffe02300007bf900001fddffff8407ffffe02300007bf900001fdd;
    assign coff[472 ] = 256'h000078c8ffffd59effff873800002a62000078c8ffffd59effff873800002a62;
    assign coff[473 ] = 256'hffffd59effff873800002a62000078c8ffffd59effff873800002a62000078c8;
    assign coff[474 ] = 256'h00003770ffff8ca1ffffc8900000735f00003770ffff8ca1ffffc8900000735f;
    assign coff[475 ] = 256'hffff8ca1ffffc8900000735f00003770ffff8ca1ffffc8900000735f00003770;
    assign coff[476 ] = 256'h00005f5effffaaa0ffffa0a20000556000005f5effffaaa0ffffa0a200005560;
    assign coff[477 ] = 256'hffffaaa0ffffa0a20000556000005f5effffaaa0ffffa0a20000556000005f5e;
    assign coff[478 ] = 256'h00000711ffff8032fffff8ef00007fce00000711ffff8032fffff8ef00007fce;
    assign coff[479 ] = 256'hffff8032fffff8ef00007fce00000711ffff8032fffff8ef00007fce00000711;
    assign coff[480 ] = 256'h00007f75fffff43cffff808b00000bc400007f75fffff43cffff808b00000bc4;
    assign coff[481 ] = 256'hfffff43cffff808b00000bc400007f75fffff43cffff808b00000bc400007f75;
    assign coff[482 ] = 256'h000051cfffff9d8effffae3100006272000051cfffff9d8effffae3100006272;
    assign coff[483 ] = 256'hffff9d8effffae3100006272000051cfffff9d8effffae3100006272000051cf;
    assign coff[484 ] = 256'h00007141ffffc45bffff8ebf00003ba500007141ffffc45bffff8ebf00003ba5;
    assign coff[485 ] = 256'hffffc45bffff8ebf00003ba500007141ffffc45bffff8ebf00003ba500007141;
    assign coff[486 ] = 256'h000025e8ffff85beffffda1800007a42000025e8ffff85beffffda1800007a42;
    assign coff[487 ] = 256'hffff85beffffda1800007a42000025e8ffff85beffffda1800007a42000025e8;
    assign coff[488 ] = 256'h00007ab7ffffdb99ffff85490000246700007ab7ffffdb99ffff854900002467;
    assign coff[489 ] = 256'hffffdb99ffff85490000246700007ab7ffffdb99ffff85490000246700007ab7;
    assign coff[490 ] = 256'h00003d08ffff8f7dffffc2f80000708300003d08ffff8f7dffffc2f800007083;
    assign coff[491 ] = 256'hffff8f7dffffc2f80000708300003d08ffff8f7dffffc2f80000708300003d08;
    assign coff[492 ] = 256'h00006371ffffaf68ffff9c8f0000509800006371ffffaf68ffff9c8f00005098;
    assign coff[493 ] = 256'hffffaf68ffff9c8f0000509800006371ffffaf68ffff9c8f0000509800006371;
    assign coff[494 ] = 256'h00000d54ffff80b2fffff2ac00007f4e00000d54ffff80b2fffff2ac00007f4e;
    assign coff[495 ] = 256'hffff80b2fffff2ac00007f4e00000d54ffff80b2fffff2ac00007f4e00000d54;
    assign coff[496 ] = 256'h00007db1ffffe7cdffff824f0000183300007db1ffffe7cdffff824f00001833;
    assign coff[497 ] = 256'hffffe7cdffff824f0000183300007db1ffffe7cdffff824f0000183300007db1;
    assign coff[498 ] = 256'h000047c4ffff9603ffffb83c000069fd000047c4ffff9603ffffb83c000069fd;
    assign coff[499 ] = 256'hffff9603ffffb83c000069fd000047c4ffff9603ffffb83c000069fd000047c4;
    assign coff[500 ] = 256'h00006addffffb98bffff95230000467500006addffffb98bffff952300004675;
    assign coff[501 ] = 256'hffffb98bffff95230000467500006addffffb98bffff95230000467500006add;
    assign coff[502 ] = 256'h000019beffff829dffffe64200007d63000019beffff829dffffe64200007d63;
    assign coff[503 ] = 256'hffff829dffffe64200007d63000019beffff829dffffe64200007d63000019be;
    assign coff[504 ] = 256'h0000768effffcfbeffff8972000030420000768effffcfbeffff897200003042;
    assign coff[505 ] = 256'hffffcfbeffff8972000030420000768effffcfbeffff8972000030420000768e;
    assign coff[506 ] = 256'h000031b5ffff8a0cffffce4b000075f4000031b5ffff8a0cffffce4b000075f4;
    assign coff[507 ] = 256'hffff8a0cffffce4b000075f4000031b5ffff8a0cffffce4b000075f4000031b5;
    assign coff[508 ] = 256'h00005b10ffffa60cffffa4f0000059f400005b10ffffa60cffffa4f0000059f4;
    assign coff[509 ] = 256'hffffa60cffffa4f0000059f400005b10ffffa60cffffa4f0000059f400005b10;
    assign coff[510 ] = 256'h000000c9ffff8001ffffff3700007fff000000c9ffff8001ffffff3700007fff;
    assign coff[511 ] = 256'hffff8001ffffff3700007fff000000c9ffff8001ffffff3700007fff000000c9;
    assign coff[512 ] = 256'h00007fffffffff9bffff80010000006500007fffffffff9bffff800100000065;
    assign coff[513 ] = 256'hffffff9bffff80010000006500007fffffffff9bffff80010000006500007fff;
    assign coff[514 ] = 256'h00005a3bffffa537ffffa5c500005ac900005a3bffffa537ffffa5c500005ac9;
    assign coff[515 ] = 256'hffffa537ffffa5c500005ac900005a3bffffa537ffffa5c500005ac900005a3b;
    assign coff[516 ] = 256'h0000761bffffcea7ffff89e5000031590000761bffffcea7ffff89e500003159;
    assign coff[517 ] = 256'hffffcea7ffff89e5000031590000761bffffcea7ffff89e5000031590000761b;
    assign coff[518 ] = 256'h0000309fffff8998ffffcf61000076680000309fffff8998ffffcf6100007668;
    assign coff[519 ] = 256'hffff8998ffffcf61000076680000309fffff8998ffffcf61000076680000309f;
    assign coff[520 ] = 256'h00007d77ffffe6a5ffff82890000195b00007d77ffffe6a5ffff82890000195b;
    assign coff[521 ] = 256'hffffe6a5ffff82890000195b00007d77ffffe6a5ffff82890000195b00007d77;
    assign coff[522 ] = 256'h000046c9ffff955bffffb93700006aa5000046c9ffff955bffffb93700006aa5;
    assign coff[523 ] = 256'hffff955bffffb93700006aa5000046c9ffff955bffffb93700006aa5000046c9;
    assign coff[524 ] = 256'h00006a36ffffb890ffff95ca0000477000006a36ffffb890ffff95ca00004770;
    assign coff[525 ] = 256'hffffb890ffff95ca0000477000006a36ffffb890ffff95ca0000477000006a36;
    assign coff[526 ] = 256'h00001896ffff8262ffffe76a00007d9e00001896ffff8262ffffe76a00007d9e;
    assign coff[527 ] = 256'hffff8262ffffe76a00007d9e00001896ffff8262ffffe76a00007d9e00001896;
    assign coff[528 ] = 256'h00007f58fffff310ffff80a800000cf000007f58fffff310ffff80a800000cf0;
    assign coff[529 ] = 256'hfffff310ffff80a800000cf000007f58fffff310ffff80a800000cf000007f58;
    assign coff[530 ] = 256'h000050e6ffff9cceffffaf1a00006332000050e6ffff9cceffffaf1a00006332;
    assign coff[531 ] = 256'hffff9cceffffaf1a00006332000050e6ffff9cceffffaf1a00006332000050e6;
    assign coff[532 ] = 256'h000070b3ffffc351ffff8f4d00003caf000070b3ffffc351ffff8f4d00003caf;
    assign coff[533 ] = 256'hffffc351ffff8f4d00003caf000070b3ffffc351ffff8f4d00003caf000070b3;
    assign coff[534 ] = 256'h000024c8ffff8566ffffdb3800007a9a000024c8ffff8566ffffdb3800007a9a;
    assign coff[535 ] = 256'hffff8566ffffdb3800007a9a000024c8ffff8566ffffdb3800007a9a000024c8;
    assign coff[536 ] = 256'h00007a60ffffda78ffff85a00000258800007a60ffffda78ffff85a000002588;
    assign coff[537 ] = 256'hffffda78ffff85a00000258800007a60ffffda78ffff85a00000258800007a60;
    assign coff[538 ] = 256'h00003bfeffff8eeeffffc4020000711200003bfeffff8eeeffffc40200007112;
    assign coff[539 ] = 256'hffff8eeeffffc4020000711200003bfeffff8eeeffffc4020000711200003bfe;
    assign coff[540 ] = 256'h000062b2ffffae7fffff9d4e00005181000062b2ffffae7fffff9d4e00005181;
    assign coff[541 ] = 256'hffffae7fffff9d4e00005181000062b2ffffae7fffff9d4e00005181000062b2;
    assign coff[542 ] = 256'h00000c28ffff8094fffff3d800007f6c00000c28ffff8094fffff3d800007f6c;
    assign coff[543 ] = 256'hffff8094fffff3d800007f6c00000c28ffff8094fffff3d800007f6c00000c28;
    assign coff[544 ] = 256'h00007fd3fffff954ffff802d000006ac00007fd3fffff954ffff802d000006ac;
    assign coff[545 ] = 256'hfffff954ffff802d000006ac00007fd3fffff954ffff802d000006ac00007fd3;
    assign coff[546 ] = 256'h000055abffffa0e5ffffaa5500005f1b000055abffffa0e5ffffaa5500005f1b;
    assign coff[547 ] = 256'hffffa0e5ffffaa5500005f1b000055abffffa0e5ffffaa5500005f1b000055ab;
    assign coff[548 ] = 256'h0000738bffffc8ebffff8c75000037150000738bffffc8ebffff8c7500003715;
    assign coff[549 ] = 256'hffffc8ebffff8c75000037150000738bffffc8ebffff8c75000037150000738b;
    assign coff[550 ] = 256'h00002ac1ffff875affffd53f000078a600002ac1ffff875affffd53f000078a6;
    assign coff[551 ] = 256'hffff875affffd53f000078a600002ac1ffff875affffd53f000078a600002ac1;
    assign coff[552 ] = 256'h00007c11ffffe085ffff83ef00001f7b00007c11ffffe085ffff83ef00001f7b;
    assign coff[553 ] = 256'hffffe085ffff83ef00001f7b00007c11ffffe085ffff83ef00001f7b00007c11;
    assign coff[554 ] = 256'h00004178ffff9202ffffbe8800006dfe00004178ffff9202ffffbe8800006dfe;
    assign coff[555 ] = 256'hffff9202ffffbe8800006dfe00004178ffff9202ffffbe8800006dfe00004178;
    assign coff[556 ] = 256'h00006693ffffb36fffff996d00004c9100006693ffffb36fffff996d00004c91;
    assign coff[557 ] = 256'hffffb36fffff996d00004c9100006693ffffb36fffff996d00004c9100006693;
    assign coff[558 ] = 256'h00001265ffff8154ffffed9b00007eac00001265ffff8154ffffed9b00007eac;
    assign coff[559 ] = 256'hffff8154ffffed9b00007eac00001265ffff8154ffffed9b00007eac00001265;
    assign coff[560 ] = 256'h00007e8effffecd5ffff81720000132b00007e8effffecd5ffff81720000132b;
    assign coff[561 ] = 256'hffffecd5ffff81720000132b00007e8effffecd5ffff81720000132b00007e8e;
    assign coff[562 ] = 256'h00004befffff98f5ffffb4110000670b00004befffff98f5ffffb4110000670b;
    assign coff[563 ] = 256'hffff98f5ffffb4110000670b00004befffff98f5ffffb4110000670b00004bef;
    assign coff[564 ] = 256'h00006d96ffffbddcffff926a0000422400006d96ffffbddcffff926a00004224;
    assign coff[565 ] = 256'hffffbddcffff926a0000422400006d96ffffbddcffff926a0000422400006d96;
    assign coff[566 ] = 256'h00001eb8ffff83beffffe14800007c4200001eb8ffff83beffffe14800007c42;
    assign coff[567 ] = 256'hffff83beffffe14800007c4200001eb8ffff83beffffe14800007c4200001eb8;
    assign coff[568 ] = 256'h00007863ffffd482ffff879d00002b7e00007863ffffd482ffff879d00002b7e;
    assign coff[569 ] = 256'hffffd482ffff879d00002b7e00007863ffffd482ffff879d00002b7e00007863;
    assign coff[570 ] = 256'h0000365fffff8c1fffffc9a1000073e10000365fffff8c1fffffc9a1000073e1;
    assign coff[571 ] = 256'hffff8c1fffffc9a1000073e10000365fffff8c1fffffc9a1000073e10000365f;
    assign coff[572 ] = 256'h00005e94ffffa9c0ffffa16c0000564000005e94ffffa9c0ffffa16c00005640;
    assign coff[573 ] = 256'hffffa9c0ffffa16c0000564000005e94ffffa9c0ffffa16c0000564000005e94;
    assign coff[574 ] = 256'h000005e3ffff8023fffffa1d00007fdd000005e3ffff8023fffffa1d00007fdd;
    assign coff[575 ] = 256'hffff8023fffffa1d00007fdd000005e3ffff8023fffffa1d00007fdd000005e3;
    assign coff[576 ] = 256'h00007ff4fffffc77ffff800c0000038900007ff4fffffc77ffff800c00000389;
    assign coff[577 ] = 256'hfffffc77ffff800c0000038900007ff4fffffc77ffff800c0000038900007ff4;
    assign coff[578 ] = 256'h000057faffffa307ffffa80600005cf9000057faffffa307ffffa80600005cf9;
    assign coff[579 ] = 256'hffffa307ffffa80600005cf9000057faffffa307ffffa80600005cf9000057fa;
    assign coff[580 ] = 256'h000074dcffffcbc5ffff8b240000343b000074dcffffcbc5ffff8b240000343b;
    assign coff[581 ] = 256'hffffcbc5ffff8b240000343b000074dcffffcbc5ffff8b240000343b000074dc;
    assign coff[582 ] = 256'h00002db3ffff8870ffffd24d0000779000002db3ffff8870ffffd24d00007790;
    assign coff[583 ] = 256'hffff8870ffffd24d0000779000002db3ffff8870ffffd24d0000779000002db3;
    assign coff[584 ] = 256'h00007cceffffe392ffff833200001c6e00007cceffffe392ffff833200001c6e;
    assign coff[585 ] = 256'hffffe392ffff833200001c6e00007cceffffe392ffff833200001c6e00007cce;
    assign coff[586 ] = 256'h00004426ffff93a6ffffbbda00006c5a00004426ffff93a6ffffbbda00006c5a;
    assign coff[587 ] = 256'hffff93a6ffffbbda00006c5a00004426ffff93a6ffffbbda00006c5a00004426;
    assign coff[588 ] = 256'h0000686dffffb5faffff979300004a060000686dffffb5faffff979300004a06;
    assign coff[589 ] = 256'hffffb5faffff979300004a060000686dffffb5faffff979300004a060000686d;
    assign coff[590 ] = 256'h0000157fffff81d1ffffea8100007e2f0000157fffff81d1ffffea8100007e2f;
    assign coff[591 ] = 256'hffff81d1ffffea8100007e2f0000157fffff81d1ffffea8100007e2f0000157f;
    assign coff[592 ] = 256'h00007efdffffeff1ffff81030000100f00007efdffffeff1ffff81030000100f;
    assign coff[593 ] = 256'hffffeff1ffff81030000100f00007efdffffeff1ffff81030000100f00007efd;
    assign coff[594 ] = 256'h00004e71ffff9adaffffb18f0000652600004e71ffff9adaffffb18f00006526;
    assign coff[595 ] = 256'hffff9adaffffb18f0000652600004e71ffff9adaffffb18f0000652600004e71;
    assign coff[596 ] = 256'h00006f2dffffc091ffff90d300003f6f00006f2dffffc091ffff90d300003f6f;
    assign coff[597 ] = 256'hffffc091ffff90d300003f6f00006f2dffffc091ffff90d300003f6f00006f2d;
    assign coff[598 ] = 256'h000021c3ffff8488ffffde3d00007b78000021c3ffff8488ffffde3d00007b78;
    assign coff[599 ] = 256'hffff8488ffffde3d00007b78000021c3ffff8488ffffde3d00007b78000021c3;
    assign coff[600 ] = 256'h0000796affffd77affff8696000028860000796affffd77affff869600002886;
    assign coff[601 ] = 256'hffffd77affff8696000028860000796affffd77affff8696000028860000796a;
    assign coff[602 ] = 256'h00003933ffff8d7effffc6cd0000728200003933ffff8d7effffc6cd00007282;
    assign coff[603 ] = 256'hffff8d7effffc6cd0000728200003933ffff8d7effffc6cd0000728200003933;
    assign coff[604 ] = 256'h000060aaffffac19ffff9f56000053e7000060aaffffac19ffff9f56000053e7;
    assign coff[605 ] = 256'hffffac19ffff9f56000053e7000060aaffffac19ffff9f56000053e7000060aa;
    assign coff[606 ] = 256'h00000906ffff8052fffff6fa00007fae00000906ffff8052fffff6fa00007fae;
    assign coff[607 ] = 256'hffff8052fffff6fa00007fae00000906ffff8052fffff6fa00007fae00000906;
    assign coff[608 ] = 256'h00007fa0fffff631ffff8060000009cf00007fa0fffff631ffff8060000009cf;
    assign coff[609 ] = 256'hfffff631ffff8060000009cf00007fa0fffff631ffff8060000009cf00007fa0;
    assign coff[610 ] = 256'h0000534fffff9ed2ffffacb10000612e0000534fffff9ed2ffffacb10000612e;
    assign coff[611 ] = 256'hffff9ed2ffffacb10000612e0000534fffff9ed2ffffacb10000612e0000534f;
    assign coff[612 ] = 256'h00007228ffffc619ffff8dd8000039e700007228ffffc619ffff8dd8000039e7;
    assign coff[613 ] = 256'hffffc619ffff8dd8000039e700007228ffffc619ffff8dd8000039e700007228;
    assign coff[614 ] = 256'h000027c7ffff8656ffffd839000079aa000027c7ffff8656ffffd839000079aa;
    assign coff[615 ] = 256'hffff8656ffffd839000079aa000027c7ffff8656ffffd839000079aa000027c7;
    assign coff[616 ] = 256'h00007b42ffffdd7cffff84be0000228400007b42ffffdd7cffff84be00002284;
    assign coff[617 ] = 256'hffffdd7cffff84be0000228400007b42ffffdd7cffff84be0000228400007b42;
    assign coff[618 ] = 256'h00003ec0ffff9070ffffc14000006f9000003ec0ffff9070ffffc14000006f90;
    assign coff[619 ] = 256'hffff9070ffffc14000006f9000003ec0ffff9070ffffc14000006f9000003ec0;
    assign coff[620 ] = 256'h000064abffffb0f1ffff9b5500004f0f000064abffffb0f1ffff9b5500004f0f;
    assign coff[621 ] = 256'hffffb0f1ffff9b5500004f0f000064abffffb0f1ffff9b5500004f0f000064ab;
    assign coff[622 ] = 256'h00000f47ffff80eafffff0b900007f1600000f47ffff80eafffff0b900007f16;
    assign coff[623 ] = 256'hffff80eafffff0b900007f1600000f47ffff80eafffff0b900007f1600000f47;
    assign coff[624 ] = 256'h00007e0cffffe9bbffff81f40000164500007e0cffffe9bbffff81f400001645;
    assign coff[625 ] = 256'hffffe9bbffff81f40000164500007e0cffffe9bbffff81f40000164500007e0c;
    assign coff[626 ] = 256'h00004962ffff9720ffffb69e000068e000004962ffff9720ffffb69e000068e0;
    assign coff[627 ] = 256'hffff9720ffffb69e000068e000004962ffff9720ffffb69e000068e000004962;
    assign coff[628 ] = 256'h00006beeffffbb30ffff9412000044d000006beeffffbb30ffff9412000044d0;
    assign coff[629 ] = 256'hffffbb30ffff9412000044d000006beeffffbb30ffff9412000044d000006bee;
    assign coff[630 ] = 256'h00001ba9ffff8306ffffe45700007cfa00001ba9ffff8306ffffe45700007cfa;
    assign coff[631 ] = 256'hffff8306ffffe45700007cfa00001ba9ffff8306ffffe45700007cfa00001ba9;
    assign coff[632 ] = 256'h00007748ffffd191ffff88b800002e6f00007748ffffd191ffff88b800002e6f;
    assign coff[633 ] = 256'hffffd191ffff88b800002e6f00007748ffffd191ffff88b800002e6f00007748;
    assign coff[634 ] = 256'h00003383ffff8ad3ffffcc7d0000752d00003383ffff8ad3ffffcc7d0000752d;
    assign coff[635 ] = 256'hffff8ad3ffffcc7d0000752d00003383ffff8ad3ffffcc7d0000752d00003383;
    assign coff[636 ] = 256'h00005c6fffffa774ffffa3910000588c00005c6fffffa774ffffa3910000588c;
    assign coff[637 ] = 256'hffffa774ffffa3910000588c00005c6fffffa774ffffa3910000588c00005c6f;
    assign coff[638 ] = 256'h000002c0ffff8008fffffd4000007ff8000002c0ffff8008fffffd4000007ff8;
    assign coff[639 ] = 256'hffff8008fffffd4000007ff8000002c0ffff8008fffffd4000007ff8000002c0;
    assign coff[640 ] = 256'h00007ffcfffffe09ffff8004000001f700007ffcfffffe09ffff8004000001f7;
    assign coff[641 ] = 256'hfffffe09ffff8004000001f700007ffcfffffe09ffff8004000001f700007ffc;
    assign coff[642 ] = 256'h0000591cffffa41dffffa6e400005be30000591cffffa41dffffa6e400005be3;
    assign coff[643 ] = 256'hffffa41dffffa6e400005be30000591cffffa41dffffa6e400005be30000591c;
    assign coff[644 ] = 256'h0000757effffcd35ffff8a82000032cb0000757effffcd35ffff8a82000032cb;
    assign coff[645 ] = 256'hffffcd35ffff8a82000032cb0000757effffcd35ffff8a82000032cb0000757e;
    assign coff[646 ] = 256'h00002f2affff8902ffffd0d6000076fe00002f2affff8902ffffd0d6000076fe;
    assign coff[647 ] = 256'hffff8902ffffd0d6000076fe00002f2affff8902ffffd0d6000076fe00002f2a;
    assign coff[648 ] = 256'h00007d25ffffe51bffff82db00001ae500007d25ffffe51bffff82db00001ae5;
    assign coff[649 ] = 256'hffffe51bffff82db00001ae500007d25ffffe51bffff82db00001ae500007d25;
    assign coff[650 ] = 256'h00004579ffff947effffba8700006b8200004579ffff947effffba8700006b82;
    assign coff[651 ] = 256'hffff947effffba8700006b8200004579ffff947effffba8700006b8200004579;
    assign coff[652 ] = 256'h00006953ffffb743ffff96ad000048bd00006953ffffb743ffff96ad000048bd;
    assign coff[653 ] = 256'hffffb743ffff96ad000048bd00006953ffffb743ffff96ad000048bd00006953;
    assign coff[654 ] = 256'h0000170bffff8217ffffe8f500007de90000170bffff8217ffffe8f500007de9;
    assign coff[655 ] = 256'hffff8217ffffe8f500007de90000170bffff8217ffffe8f500007de90000170b;
    assign coff[656 ] = 256'h00007f2dfffff180ffff80d300000e8000007f2dfffff180ffff80d300000e80;
    assign coff[657 ] = 256'hfffff180ffff80d300000e8000007f2dfffff180ffff80d300000e8000007f2d;
    assign coff[658 ] = 256'h00004fadffff9bd2ffffb0530000642e00004fadffff9bd2ffffb0530000642e;
    assign coff[659 ] = 256'hffff9bd2ffffb0530000642e00004fadffff9bd2ffffb0530000642e00004fad;
    assign coff[660 ] = 256'h00006ff2ffffc1f0ffff900e00003e1000006ff2ffffc1f0ffff900e00003e10;
    assign coff[661 ] = 256'hffffc1f0ffff900e00003e1000006ff2ffffc1f0ffff900e00003e1000006ff2;
    assign coff[662 ] = 256'h00002346ffff84f5ffffdcba00007b0b00002346ffff84f5ffffdcba00007b0b;
    assign coff[663 ] = 256'hffff84f5ffffdcba00007b0b00002346ffff84f5ffffdcba00007b0b00002346;
    assign coff[664 ] = 256'h000079e7ffffd8f8ffff861900002708000079e7ffffd8f8ffff861900002708;
    assign coff[665 ] = 256'hffffd8f8ffff861900002708000079e7ffffd8f8ffff861900002708000079e7;
    assign coff[666 ] = 256'h00003a9affff8e34ffffc566000071cc00003a9affff8e34ffffc566000071cc;
    assign coff[667 ] = 256'hffff8e34ffffc566000071cc00003a9affff8e34ffffc566000071cc00003a9a;
    assign coff[668 ] = 256'h000061b0ffffad4affff9e50000052b6000061b0ffffad4affff9e50000052b6;
    assign coff[669 ] = 256'hffffad4affff9e50000052b6000061b0ffffad4affff9e50000052b6000061b0;
    assign coff[670 ] = 256'h00000a97ffff8070fffff56900007f9000000a97ffff8070fffff56900007f90;
    assign coff[671 ] = 256'hffff8070fffff56900007f9000000a97ffff8070fffff56900007f9000000a97;
    assign coff[672 ] = 256'h00007fbcfffff7c2ffff80440000083e00007fbcfffff7c2ffff80440000083e;
    assign coff[673 ] = 256'hfffff7c2ffff80440000083e00007fbcfffff7c2ffff80440000083e00007fbc;
    assign coff[674 ] = 256'h0000547fffff9fdaffffab81000060260000547fffff9fdaffffab8100006026;
    assign coff[675 ] = 256'hffff9fdaffffab81000060260000547fffff9fdaffffab81000060260000547f;
    assign coff[676 ] = 256'h000072dcffffc781ffff8d240000387f000072dcffffc781ffff8d240000387f;
    assign coff[677 ] = 256'hffffc781ffff8d240000387f000072dcffffc781ffff8d240000387f000072dc;
    assign coff[678 ] = 256'h00002945ffff86d6ffffd6bb0000792a00002945ffff86d6ffffd6bb0000792a;
    assign coff[679 ] = 256'hffff86d6ffffd6bb0000792a00002945ffff86d6ffffd6bb0000792a00002945;
    assign coff[680 ] = 256'h00007bacffffdeffffff84540000210100007bacffffdeffffff845400002101;
    assign coff[681 ] = 256'hffffdeffffff84540000210100007bacffffdeffffff84540000210100007bac;
    assign coff[682 ] = 256'h0000401dffff9137ffffbfe300006ec90000401dffff9137ffffbfe300006ec9;
    assign coff[683 ] = 256'hffff9137ffffbfe300006ec90000401dffff9137ffffbfe300006ec90000401d;
    assign coff[684 ] = 256'h000065a1ffffb22fffff9a5f00004dd1000065a1ffffb22fffff9a5f00004dd1;
    assign coff[685 ] = 256'hffffb22fffff9a5f00004dd1000065a1ffffb22fffff9a5f00004dd1000065a1;
    assign coff[686 ] = 256'h000010d6ffff811dffffef2a00007ee3000010d6ffff811dffffef2a00007ee3;
    assign coff[687 ] = 256'hffff811dffffef2a00007ee3000010d6ffff811dffffef2a00007ee3000010d6;
    assign coff[688 ] = 256'h00007e50ffffeb47ffff81b0000014b900007e50ffffeb47ffff81b0000014b9;
    assign coff[689 ] = 256'hffffeb47ffff81b0000014b900007e50ffffeb47ffff81b0000014b900007e50;
    assign coff[690 ] = 256'h00004aaaffff9808ffffb556000067f800004aaaffff9808ffffb556000067f8;
    assign coff[691 ] = 256'hffff9808ffffb556000067f800004aaaffff9808ffffb556000067f800004aaa;
    assign coff[692 ] = 256'h00006cc4ffffbc85ffff933c0000437b00006cc4ffffbc85ffff933c0000437b;
    assign coff[693 ] = 256'hffffbc85ffff933c0000437b00006cc4ffffbc85ffff933c0000437b00006cc4;
    assign coff[694 ] = 256'h00001d31ffff8360ffffe2cf00007ca000001d31ffff8360ffffe2cf00007ca0;
    assign coff[695 ] = 256'hffff8360ffffe2cf00007ca000001d31ffff8360ffffe2cf00007ca000001d31;
    assign coff[696 ] = 256'h000077d8ffffd309ffff882800002cf7000077d8ffffd309ffff882800002cf7;
    assign coff[697 ] = 256'hffffd309ffff882800002cf7000077d8ffffd309ffff882800002cf7000077d8;
    assign coff[698 ] = 256'h000034f2ffff8b77ffffcb0e00007489000034f2ffff8b77ffffcb0e00007489;
    assign coff[699 ] = 256'hffff8b77ffffcb0e00007489000034f2ffff8b77ffffcb0e00007489000034f2;
    assign coff[700 ] = 256'h00005d83ffffa899ffffa27d0000576700005d83ffffa899ffffa27d00005767;
    assign coff[701 ] = 256'hffffa899ffffa27d0000576700005d83ffffa899ffffa27d0000576700005d83;
    assign coff[702 ] = 256'h00000452ffff8013fffffbae00007fed00000452ffff8013fffffbae00007fed;
    assign coff[703 ] = 256'hffff8013fffffbae00007fed00000452ffff8013fffffbae00007fed00000452;
    assign coff[704 ] = 256'h00007fe6fffffae5ffff801a0000051b00007fe6fffffae5ffff801a0000051b;
    assign coff[705 ] = 256'hfffffae5ffff801a0000051b00007fe6fffffae5ffff801a0000051b00007fe6;
    assign coff[706 ] = 256'h000056d4ffffa1f4ffffa92c00005e0c000056d4ffffa1f4ffffa92c00005e0c;
    assign coff[707 ] = 256'hffffa1f4ffffa92c00005e0c000056d4ffffa1f4ffffa92c00005e0c000056d4;
    assign coff[708 ] = 256'h00007436ffffca57ffff8bca000035a900007436ffffca57ffff8bca000035a9;
    assign coff[709 ] = 256'hffffca57ffff8bca000035a900007436ffffca57ffff8bca000035a900007436;
    assign coff[710 ] = 256'h00002c3bffff87e2ffffd3c50000781e00002c3bffff87e2ffffd3c50000781e;
    assign coff[711 ] = 256'hffff87e2ffffd3c50000781e00002c3bffff87e2ffffd3c50000781e00002c3b;
    assign coff[712 ] = 256'h00007c72ffffe20bffff838e00001df500007c72ffffe20bffff838e00001df5;
    assign coff[713 ] = 256'hffffe20bffff838e00001df500007c72ffffe20bffff838e00001df500007c72;
    assign coff[714 ] = 256'h000042d0ffff92d2ffffbd3000006d2e000042d0ffff92d2ffffbd3000006d2e;
    assign coff[715 ] = 256'hffff92d2ffffbd3000006d2e000042d0ffff92d2ffffbd3000006d2e000042d0;
    assign coff[716 ] = 256'h00006782ffffb4b3ffff987e00004b4d00006782ffffb4b3ffff987e00004b4d;
    assign coff[717 ] = 256'hffffb4b3ffff987e00004b4d00006782ffffb4b3ffff987e00004b4d00006782;
    assign coff[718 ] = 256'h000013f2ffff8190ffffec0e00007e70000013f2ffff8190ffffec0e00007e70;
    assign coff[719 ] = 256'hffff8190ffffec0e00007e70000013f2ffff8190ffffec0e00007e70000013f2;
    assign coff[720 ] = 256'h00007ec8ffffee62ffff81380000119e00007ec8ffffee62ffff81380000119e;
    assign coff[721 ] = 256'hffffee62ffff81380000119e00007ec8ffffee62ffff81380000119e00007ec8;
    assign coff[722 ] = 256'h00004d31ffff99e5ffffb2cf0000661b00004d31ffff99e5ffffb2cf0000661b;
    assign coff[723 ] = 256'hffff99e5ffffb2cf0000661b00004d31ffff99e5ffffb2cf0000661b00004d31;
    assign coff[724 ] = 256'h00006e64ffffbf35ffff919c000040cb00006e64ffffbf35ffff919c000040cb;
    assign coff[725 ] = 256'hffffbf35ffff919c000040cb00006e64ffffbf35ffff919c000040cb00006e64;
    assign coff[726 ] = 256'h0000203effff8421ffffdfc200007bdf0000203effff8421ffffdfc200007bdf;
    assign coff[727 ] = 256'hffff8421ffffdfc200007bdf0000203effff8421ffffdfc200007bdf0000203e;
    assign coff[728 ] = 256'h000078e9ffffd5fdffff871700002a03000078e9ffffd5fdffff871700002a03;
    assign coff[729 ] = 256'hffffd5fdffff871700002a03000078e9ffffd5fdffff871700002a03000078e9;
    assign coff[730 ] = 256'h000037caffff8cccffffc83600007334000037caffff8cccffffc83600007334;
    assign coff[731 ] = 256'hffff8cccffffc83600007334000037caffff8cccffffc83600007334000037ca;
    assign coff[732 ] = 256'h00005fa1ffffaaebffffa05f0000551500005fa1ffffaaebffffa05f00005515;
    assign coff[733 ] = 256'hffffaaebffffa05f0000551500005fa1ffffaaebffffa05f0000551500005fa1;
    assign coff[734 ] = 256'h00000775ffff8038fffff88b00007fc800000775ffff8038fffff88b00007fc8;
    assign coff[735 ] = 256'hffff8038fffff88b00007fc800000775ffff8038fffff88b00007fc800000775;
    assign coff[736 ] = 256'h00007f7efffff4a0ffff808200000b6000007f7efffff4a0ffff808200000b60;
    assign coff[737 ] = 256'hfffff4a0ffff808200000b6000007f7efffff4a0ffff808200000b6000007f7e;
    assign coff[738 ] = 256'h0000521cffff9dceffffade4000062320000521cffff9dceffffade400006232;
    assign coff[739 ] = 256'hffff9dceffffade4000062320000521cffff9dceffffade4000062320000521c;
    assign coff[740 ] = 256'h00007170ffffc4b4ffff8e9000003b4c00007170ffffc4b4ffff8e9000003b4c;
    assign coff[741 ] = 256'hffffc4b4ffff8e9000003b4c00007170ffffc4b4ffff8e9000003b4c00007170;
    assign coff[742 ] = 256'h00002648ffff85dcffffd9b800007a2400002648ffff85dcffffd9b800007a24;
    assign coff[743 ] = 256'hffff85dcffffd9b800007a2400002648ffff85dcffffd9b800007a2400002648;
    assign coff[744 ] = 256'h00007ad3ffffdbf9ffff852d0000240700007ad3ffffdbf9ffff852d00002407;
    assign coff[745 ] = 256'hffffdbf9ffff852d0000240700007ad3ffffdbf9ffff852d0000240700007ad3;
    assign coff[746 ] = 256'h00003d60ffff8fadffffc2a00000705300003d60ffff8fadffffc2a000007053;
    assign coff[747 ] = 256'hffff8fadffffc2a00000705300003d60ffff8fadffffc2a00000705300003d60;
    assign coff[748 ] = 256'h000063b0ffffafb6ffff9c500000504a000063b0ffffafb6ffff9c500000504a;
    assign coff[749 ] = 256'hffffafb6ffff9c500000504a000063b0ffffafb6ffff9c500000504a000063b0;
    assign coff[750 ] = 256'h00000db8ffff80bdfffff24800007f4300000db8ffff80bdfffff24800007f43;
    assign coff[751 ] = 256'hffff80bdfffff24800007f4300000db8ffff80bdfffff24800007f4300000db8;
    assign coff[752 ] = 256'h00007dc4ffffe82fffff823c000017d100007dc4ffffe82fffff823c000017d1;
    assign coff[753 ] = 256'hffffe82fffff823c000017d100007dc4ffffe82fffff823c000017d100007dc4;
    assign coff[754 ] = 256'h00004817ffff963bffffb7e9000069c500004817ffff963bffffb7e9000069c5;
    assign coff[755 ] = 256'hffff963bffffb7e9000069c500004817ffff963bffffb7e9000069c500004817;
    assign coff[756 ] = 256'h00006b14ffffb9dfffff94ec0000462100006b14ffffb9dfffff94ec00004621;
    assign coff[757 ] = 256'hffffb9dfffff94ec0000462100006b14ffffb9dfffff94ec0000462100006b14;
    assign coff[758 ] = 256'h00001a20ffff82b2ffffe5e000007d4e00001a20ffff82b2ffffe5e000007d4e;
    assign coff[759 ] = 256'hffff82b2ffffe5e000007d4e00001a20ffff82b2ffffe5e000007d4e00001a20;
    assign coff[760 ] = 256'h000076b4ffffd01bffff894c00002fe5000076b4ffffd01bffff894c00002fe5;
    assign coff[761 ] = 256'hffffd01bffff894c00002fe5000076b4ffffd01bffff894c00002fe5000076b4;
    assign coff[762 ] = 256'h00003212ffff8a33ffffcdee000075cd00003212ffff8a33ffffcdee000075cd;
    assign coff[763 ] = 256'hffff8a33ffffcdee000075cd00003212ffff8a33ffffcdee000075cd00003212;
    assign coff[764 ] = 256'h00005b57ffffa654ffffa4a9000059ac00005b57ffffa654ffffa4a9000059ac;
    assign coff[765 ] = 256'hffffa654ffffa4a9000059ac00005b57ffffa654ffffa4a9000059ac00005b57;
    assign coff[766 ] = 256'h0000012effff8001fffffed200007fff0000012effff8001fffffed200007fff;
    assign coff[767 ] = 256'hffff8001fffffed200007fff0000012effff8001fffffed200007fff0000012e;
    assign coff[768 ] = 256'h00007ffffffffed2ffff80010000012e00007ffffffffed2ffff80010000012e;
    assign coff[769 ] = 256'hfffffed2ffff80010000012e00007ffffffffed2ffff80010000012e00007fff;
    assign coff[770 ] = 256'h000059acffffa4a9ffffa65400005b57000059acffffa4a9ffffa65400005b57;
    assign coff[771 ] = 256'hffffa4a9ffffa65400005b57000059acffffa4a9ffffa65400005b57000059ac;
    assign coff[772 ] = 256'h000075cdffffcdeeffff8a3300003212000075cdffffcdeeffff8a3300003212;
    assign coff[773 ] = 256'hffffcdeeffff8a3300003212000075cdffffcdeeffff8a3300003212000075cd;
    assign coff[774 ] = 256'h00002fe5ffff894cffffd01b000076b400002fe5ffff894cffffd01b000076b4;
    assign coff[775 ] = 256'hffff894cffffd01b000076b400002fe5ffff894cffffd01b000076b400002fe5;
    assign coff[776 ] = 256'h00007d4effffe5e0ffff82b200001a2000007d4effffe5e0ffff82b200001a20;
    assign coff[777 ] = 256'hffffe5e0ffff82b200001a2000007d4effffe5e0ffff82b200001a2000007d4e;
    assign coff[778 ] = 256'h00004621ffff94ecffffb9df00006b1400004621ffff94ecffffb9df00006b14;
    assign coff[779 ] = 256'hffff94ecffffb9df00006b1400004621ffff94ecffffb9df00006b1400004621;
    assign coff[780 ] = 256'h000069c5ffffb7e9ffff963b00004817000069c5ffffb7e9ffff963b00004817;
    assign coff[781 ] = 256'hffffb7e9ffff963b00004817000069c5ffffb7e9ffff963b00004817000069c5;
    assign coff[782 ] = 256'h000017d1ffff823cffffe82f00007dc4000017d1ffff823cffffe82f00007dc4;
    assign coff[783 ] = 256'hffff823cffffe82f00007dc4000017d1ffff823cffffe82f00007dc4000017d1;
    assign coff[784 ] = 256'h00007f43fffff248ffff80bd00000db800007f43fffff248ffff80bd00000db8;
    assign coff[785 ] = 256'hfffff248ffff80bd00000db800007f43fffff248ffff80bd00000db800007f43;
    assign coff[786 ] = 256'h0000504affff9c50ffffafb6000063b00000504affff9c50ffffafb6000063b0;
    assign coff[787 ] = 256'hffff9c50ffffafb6000063b00000504affff9c50ffffafb6000063b00000504a;
    assign coff[788 ] = 256'h00007053ffffc2a0ffff8fad00003d6000007053ffffc2a0ffff8fad00003d60;
    assign coff[789 ] = 256'hffffc2a0ffff8fad00003d6000007053ffffc2a0ffff8fad00003d6000007053;
    assign coff[790 ] = 256'h00002407ffff852dffffdbf900007ad300002407ffff852dffffdbf900007ad3;
    assign coff[791 ] = 256'hffff852dffffdbf900007ad300002407ffff852dffffdbf900007ad300002407;
    assign coff[792 ] = 256'h00007a24ffffd9b8ffff85dc0000264800007a24ffffd9b8ffff85dc00002648;
    assign coff[793 ] = 256'hffffd9b8ffff85dc0000264800007a24ffffd9b8ffff85dc0000264800007a24;
    assign coff[794 ] = 256'h00003b4cffff8e90ffffc4b40000717000003b4cffff8e90ffffc4b400007170;
    assign coff[795 ] = 256'hffff8e90ffffc4b40000717000003b4cffff8e90ffffc4b40000717000003b4c;
    assign coff[796 ] = 256'h00006232ffffade4ffff9dce0000521c00006232ffffade4ffff9dce0000521c;
    assign coff[797 ] = 256'hffffade4ffff9dce0000521c00006232ffffade4ffff9dce0000521c00006232;
    assign coff[798 ] = 256'h00000b60ffff8082fffff4a000007f7e00000b60ffff8082fffff4a000007f7e;
    assign coff[799 ] = 256'hffff8082fffff4a000007f7e00000b60ffff8082fffff4a000007f7e00000b60;
    assign coff[800 ] = 256'h00007fc8fffff88bffff80380000077500007fc8fffff88bffff803800000775;
    assign coff[801 ] = 256'hfffff88bffff80380000077500007fc8fffff88bffff80380000077500007fc8;
    assign coff[802 ] = 256'h00005515ffffa05fffffaaeb00005fa100005515ffffa05fffffaaeb00005fa1;
    assign coff[803 ] = 256'hffffa05fffffaaeb00005fa100005515ffffa05fffffaaeb00005fa100005515;
    assign coff[804 ] = 256'h00007334ffffc836ffff8ccc000037ca00007334ffffc836ffff8ccc000037ca;
    assign coff[805 ] = 256'hffffc836ffff8ccc000037ca00007334ffffc836ffff8ccc000037ca00007334;
    assign coff[806 ] = 256'h00002a03ffff8717ffffd5fd000078e900002a03ffff8717ffffd5fd000078e9;
    assign coff[807 ] = 256'hffff8717ffffd5fd000078e900002a03ffff8717ffffd5fd000078e900002a03;
    assign coff[808 ] = 256'h00007bdfffffdfc2ffff84210000203e00007bdfffffdfc2ffff84210000203e;
    assign coff[809 ] = 256'hffffdfc2ffff84210000203e00007bdfffffdfc2ffff84210000203e00007bdf;
    assign coff[810 ] = 256'h000040cbffff919cffffbf3500006e64000040cbffff919cffffbf3500006e64;
    assign coff[811 ] = 256'hffff919cffffbf3500006e64000040cbffff919cffffbf3500006e64000040cb;
    assign coff[812 ] = 256'h0000661bffffb2cfffff99e500004d310000661bffffb2cfffff99e500004d31;
    assign coff[813 ] = 256'hffffb2cfffff99e500004d310000661bffffb2cfffff99e500004d310000661b;
    assign coff[814 ] = 256'h0000119effff8138ffffee6200007ec80000119effff8138ffffee6200007ec8;
    assign coff[815 ] = 256'hffff8138ffffee6200007ec80000119effff8138ffffee6200007ec80000119e;
    assign coff[816 ] = 256'h00007e70ffffec0effff8190000013f200007e70ffffec0effff8190000013f2;
    assign coff[817 ] = 256'hffffec0effff8190000013f200007e70ffffec0effff8190000013f200007e70;
    assign coff[818 ] = 256'h00004b4dffff987effffb4b30000678200004b4dffff987effffb4b300006782;
    assign coff[819 ] = 256'hffff987effffb4b30000678200004b4dffff987effffb4b30000678200004b4d;
    assign coff[820 ] = 256'h00006d2effffbd30ffff92d2000042d000006d2effffbd30ffff92d2000042d0;
    assign coff[821 ] = 256'hffffbd30ffff92d2000042d000006d2effffbd30ffff92d2000042d000006d2e;
    assign coff[822 ] = 256'h00001df5ffff838effffe20b00007c7200001df5ffff838effffe20b00007c72;
    assign coff[823 ] = 256'hffff838effffe20b00007c7200001df5ffff838effffe20b00007c7200001df5;
    assign coff[824 ] = 256'h0000781effffd3c5ffff87e200002c3b0000781effffd3c5ffff87e200002c3b;
    assign coff[825 ] = 256'hffffd3c5ffff87e200002c3b0000781effffd3c5ffff87e200002c3b0000781e;
    assign coff[826 ] = 256'h000035a9ffff8bcaffffca5700007436000035a9ffff8bcaffffca5700007436;
    assign coff[827 ] = 256'hffff8bcaffffca5700007436000035a9ffff8bcaffffca5700007436000035a9;
    assign coff[828 ] = 256'h00005e0cffffa92cffffa1f4000056d400005e0cffffa92cffffa1f4000056d4;
    assign coff[829 ] = 256'hffffa92cffffa1f4000056d400005e0cffffa92cffffa1f4000056d400005e0c;
    assign coff[830 ] = 256'h0000051bffff801afffffae500007fe60000051bffff801afffffae500007fe6;
    assign coff[831 ] = 256'hffff801afffffae500007fe60000051bffff801afffffae500007fe60000051b;
    assign coff[832 ] = 256'h00007fedfffffbaeffff80130000045200007fedfffffbaeffff801300000452;
    assign coff[833 ] = 256'hfffffbaeffff80130000045200007fedfffffbaeffff80130000045200007fed;
    assign coff[834 ] = 256'h00005767ffffa27dffffa89900005d8300005767ffffa27dffffa89900005d83;
    assign coff[835 ] = 256'hffffa27dffffa89900005d8300005767ffffa27dffffa89900005d8300005767;
    assign coff[836 ] = 256'h00007489ffffcb0effff8b77000034f200007489ffffcb0effff8b77000034f2;
    assign coff[837 ] = 256'hffffcb0effff8b77000034f200007489ffffcb0effff8b77000034f200007489;
    assign coff[838 ] = 256'h00002cf7ffff8828ffffd309000077d800002cf7ffff8828ffffd309000077d8;
    assign coff[839 ] = 256'hffff8828ffffd309000077d800002cf7ffff8828ffffd309000077d800002cf7;
    assign coff[840 ] = 256'h00007ca0ffffe2cfffff836000001d3100007ca0ffffe2cfffff836000001d31;
    assign coff[841 ] = 256'hffffe2cfffff836000001d3100007ca0ffffe2cfffff836000001d3100007ca0;
    assign coff[842 ] = 256'h0000437bffff933cffffbc8500006cc40000437bffff933cffffbc8500006cc4;
    assign coff[843 ] = 256'hffff933cffffbc8500006cc40000437bffff933cffffbc8500006cc40000437b;
    assign coff[844 ] = 256'h000067f8ffffb556ffff980800004aaa000067f8ffffb556ffff980800004aaa;
    assign coff[845 ] = 256'hffffb556ffff980800004aaa000067f8ffffb556ffff980800004aaa000067f8;
    assign coff[846 ] = 256'h000014b9ffff81b0ffffeb4700007e50000014b9ffff81b0ffffeb4700007e50;
    assign coff[847 ] = 256'hffff81b0ffffeb4700007e50000014b9ffff81b0ffffeb4700007e50000014b9;
    assign coff[848 ] = 256'h00007ee3ffffef2affff811d000010d600007ee3ffffef2affff811d000010d6;
    assign coff[849 ] = 256'hffffef2affff811d000010d600007ee3ffffef2affff811d000010d600007ee3;
    assign coff[850 ] = 256'h00004dd1ffff9a5fffffb22f000065a100004dd1ffff9a5fffffb22f000065a1;
    assign coff[851 ] = 256'hffff9a5fffffb22f000065a100004dd1ffff9a5fffffb22f000065a100004dd1;
    assign coff[852 ] = 256'h00006ec9ffffbfe3ffff91370000401d00006ec9ffffbfe3ffff91370000401d;
    assign coff[853 ] = 256'hffffbfe3ffff91370000401d00006ec9ffffbfe3ffff91370000401d00006ec9;
    assign coff[854 ] = 256'h00002101ffff8454ffffdeff00007bac00002101ffff8454ffffdeff00007bac;
    assign coff[855 ] = 256'hffff8454ffffdeff00007bac00002101ffff8454ffffdeff00007bac00002101;
    assign coff[856 ] = 256'h0000792affffd6bbffff86d6000029450000792affffd6bbffff86d600002945;
    assign coff[857 ] = 256'hffffd6bbffff86d6000029450000792affffd6bbffff86d6000029450000792a;
    assign coff[858 ] = 256'h0000387fffff8d24ffffc781000072dc0000387fffff8d24ffffc781000072dc;
    assign coff[859 ] = 256'hffff8d24ffffc781000072dc0000387fffff8d24ffffc781000072dc0000387f;
    assign coff[860 ] = 256'h00006026ffffab81ffff9fda0000547f00006026ffffab81ffff9fda0000547f;
    assign coff[861 ] = 256'hffffab81ffff9fda0000547f00006026ffffab81ffff9fda0000547f00006026;
    assign coff[862 ] = 256'h0000083effff8044fffff7c200007fbc0000083effff8044fffff7c200007fbc;
    assign coff[863 ] = 256'hffff8044fffff7c200007fbc0000083effff8044fffff7c200007fbc0000083e;
    assign coff[864 ] = 256'h00007f90fffff569ffff807000000a9700007f90fffff569ffff807000000a97;
    assign coff[865 ] = 256'hfffff569ffff807000000a9700007f90fffff569ffff807000000a9700007f90;
    assign coff[866 ] = 256'h000052b6ffff9e50ffffad4a000061b0000052b6ffff9e50ffffad4a000061b0;
    assign coff[867 ] = 256'hffff9e50ffffad4a000061b0000052b6ffff9e50ffffad4a000061b0000052b6;
    assign coff[868 ] = 256'h000071ccffffc566ffff8e3400003a9a000071ccffffc566ffff8e3400003a9a;
    assign coff[869 ] = 256'hffffc566ffff8e3400003a9a000071ccffffc566ffff8e3400003a9a000071cc;
    assign coff[870 ] = 256'h00002708ffff8619ffffd8f8000079e700002708ffff8619ffffd8f8000079e7;
    assign coff[871 ] = 256'hffff8619ffffd8f8000079e700002708ffff8619ffffd8f8000079e700002708;
    assign coff[872 ] = 256'h00007b0bffffdcbaffff84f50000234600007b0bffffdcbaffff84f500002346;
    assign coff[873 ] = 256'hffffdcbaffff84f50000234600007b0bffffdcbaffff84f50000234600007b0b;
    assign coff[874 ] = 256'h00003e10ffff900effffc1f000006ff200003e10ffff900effffc1f000006ff2;
    assign coff[875 ] = 256'hffff900effffc1f000006ff200003e10ffff900effffc1f000006ff200003e10;
    assign coff[876 ] = 256'h0000642effffb053ffff9bd200004fad0000642effffb053ffff9bd200004fad;
    assign coff[877 ] = 256'hffffb053ffff9bd200004fad0000642effffb053ffff9bd200004fad0000642e;
    assign coff[878 ] = 256'h00000e80ffff80d3fffff18000007f2d00000e80ffff80d3fffff18000007f2d;
    assign coff[879 ] = 256'hffff80d3fffff18000007f2d00000e80ffff80d3fffff18000007f2d00000e80;
    assign coff[880 ] = 256'h00007de9ffffe8f5ffff82170000170b00007de9ffffe8f5ffff82170000170b;
    assign coff[881 ] = 256'hffffe8f5ffff82170000170b00007de9ffffe8f5ffff82170000170b00007de9;
    assign coff[882 ] = 256'h000048bdffff96adffffb74300006953000048bdffff96adffffb74300006953;
    assign coff[883 ] = 256'hffff96adffffb74300006953000048bdffff96adffffb74300006953000048bd;
    assign coff[884 ] = 256'h00006b82ffffba87ffff947e0000457900006b82ffffba87ffff947e00004579;
    assign coff[885 ] = 256'hffffba87ffff947e0000457900006b82ffffba87ffff947e0000457900006b82;
    assign coff[886 ] = 256'h00001ae5ffff82dbffffe51b00007d2500001ae5ffff82dbffffe51b00007d25;
    assign coff[887 ] = 256'hffff82dbffffe51b00007d2500001ae5ffff82dbffffe51b00007d2500001ae5;
    assign coff[888 ] = 256'h000076feffffd0d6ffff890200002f2a000076feffffd0d6ffff890200002f2a;
    assign coff[889 ] = 256'hffffd0d6ffff890200002f2a000076feffffd0d6ffff890200002f2a000076fe;
    assign coff[890 ] = 256'h000032cbffff8a82ffffcd350000757e000032cbffff8a82ffffcd350000757e;
    assign coff[891 ] = 256'hffff8a82ffffcd350000757e000032cbffff8a82ffffcd350000757e000032cb;
    assign coff[892 ] = 256'h00005be3ffffa6e4ffffa41d0000591c00005be3ffffa6e4ffffa41d0000591c;
    assign coff[893 ] = 256'hffffa6e4ffffa41d0000591c00005be3ffffa6e4ffffa41d0000591c00005be3;
    assign coff[894 ] = 256'h000001f7ffff8004fffffe0900007ffc000001f7ffff8004fffffe0900007ffc;
    assign coff[895 ] = 256'hffff8004fffffe0900007ffc000001f7ffff8004fffffe0900007ffc000001f7;
    assign coff[896 ] = 256'h00007ff8fffffd40ffff8008000002c000007ff8fffffd40ffff8008000002c0;
    assign coff[897 ] = 256'hfffffd40ffff8008000002c000007ff8fffffd40ffff8008000002c000007ff8;
    assign coff[898 ] = 256'h0000588cffffa391ffffa77400005c6f0000588cffffa391ffffa77400005c6f;
    assign coff[899 ] = 256'hffffa391ffffa77400005c6f0000588cffffa391ffffa77400005c6f0000588c;
    assign coff[900 ] = 256'h0000752dffffcc7dffff8ad3000033830000752dffffcc7dffff8ad300003383;
    assign coff[901 ] = 256'hffffcc7dffff8ad3000033830000752dffffcc7dffff8ad3000033830000752d;
    assign coff[902 ] = 256'h00002e6fffff88b8ffffd1910000774800002e6fffff88b8ffffd19100007748;
    assign coff[903 ] = 256'hffff88b8ffffd1910000774800002e6fffff88b8ffffd1910000774800002e6f;
    assign coff[904 ] = 256'h00007cfaffffe457ffff830600001ba900007cfaffffe457ffff830600001ba9;
    assign coff[905 ] = 256'hffffe457ffff830600001ba900007cfaffffe457ffff830600001ba900007cfa;
    assign coff[906 ] = 256'h000044d0ffff9412ffffbb3000006bee000044d0ffff9412ffffbb3000006bee;
    assign coff[907 ] = 256'hffff9412ffffbb3000006bee000044d0ffff9412ffffbb3000006bee000044d0;
    assign coff[908 ] = 256'h000068e0ffffb69effff972000004962000068e0ffffb69effff972000004962;
    assign coff[909 ] = 256'hffffb69effff972000004962000068e0ffffb69effff972000004962000068e0;
    assign coff[910 ] = 256'h00001645ffff81f4ffffe9bb00007e0c00001645ffff81f4ffffe9bb00007e0c;
    assign coff[911 ] = 256'hffff81f4ffffe9bb00007e0c00001645ffff81f4ffffe9bb00007e0c00001645;
    assign coff[912 ] = 256'h00007f16fffff0b9ffff80ea00000f4700007f16fffff0b9ffff80ea00000f47;
    assign coff[913 ] = 256'hfffff0b9ffff80ea00000f4700007f16fffff0b9ffff80ea00000f4700007f16;
    assign coff[914 ] = 256'h00004f0fffff9b55ffffb0f1000064ab00004f0fffff9b55ffffb0f1000064ab;
    assign coff[915 ] = 256'hffff9b55ffffb0f1000064ab00004f0fffff9b55ffffb0f1000064ab00004f0f;
    assign coff[916 ] = 256'h00006f90ffffc140ffff907000003ec000006f90ffffc140ffff907000003ec0;
    assign coff[917 ] = 256'hffffc140ffff907000003ec000006f90ffffc140ffff907000003ec000006f90;
    assign coff[918 ] = 256'h00002284ffff84beffffdd7c00007b4200002284ffff84beffffdd7c00007b42;
    assign coff[919 ] = 256'hffff84beffffdd7c00007b4200002284ffff84beffffdd7c00007b4200002284;
    assign coff[920 ] = 256'h000079aaffffd839ffff8656000027c7000079aaffffd839ffff8656000027c7;
    assign coff[921 ] = 256'hffffd839ffff8656000027c7000079aaffffd839ffff8656000027c7000079aa;
    assign coff[922 ] = 256'h000039e7ffff8dd8ffffc61900007228000039e7ffff8dd8ffffc61900007228;
    assign coff[923 ] = 256'hffff8dd8ffffc61900007228000039e7ffff8dd8ffffc61900007228000039e7;
    assign coff[924 ] = 256'h0000612effffacb1ffff9ed20000534f0000612effffacb1ffff9ed20000534f;
    assign coff[925 ] = 256'hffffacb1ffff9ed20000534f0000612effffacb1ffff9ed20000534f0000612e;
    assign coff[926 ] = 256'h000009cfffff8060fffff63100007fa0000009cfffff8060fffff63100007fa0;
    assign coff[927 ] = 256'hffff8060fffff63100007fa0000009cfffff8060fffff63100007fa0000009cf;
    assign coff[928 ] = 256'h00007faefffff6faffff80520000090600007faefffff6faffff805200000906;
    assign coff[929 ] = 256'hfffff6faffff80520000090600007faefffff6faffff80520000090600007fae;
    assign coff[930 ] = 256'h000053e7ffff9f56ffffac19000060aa000053e7ffff9f56ffffac19000060aa;
    assign coff[931 ] = 256'hffff9f56ffffac19000060aa000053e7ffff9f56ffffac19000060aa000053e7;
    assign coff[932 ] = 256'h00007282ffffc6cdffff8d7e0000393300007282ffffc6cdffff8d7e00003933;
    assign coff[933 ] = 256'hffffc6cdffff8d7e0000393300007282ffffc6cdffff8d7e0000393300007282;
    assign coff[934 ] = 256'h00002886ffff8696ffffd77a0000796a00002886ffff8696ffffd77a0000796a;
    assign coff[935 ] = 256'hffff8696ffffd77a0000796a00002886ffff8696ffffd77a0000796a00002886;
    assign coff[936 ] = 256'h00007b78ffffde3dffff8488000021c300007b78ffffde3dffff8488000021c3;
    assign coff[937 ] = 256'hffffde3dffff8488000021c300007b78ffffde3dffff8488000021c300007b78;
    assign coff[938 ] = 256'h00003f6fffff90d3ffffc09100006f2d00003f6fffff90d3ffffc09100006f2d;
    assign coff[939 ] = 256'hffff90d3ffffc09100006f2d00003f6fffff90d3ffffc09100006f2d00003f6f;
    assign coff[940 ] = 256'h00006526ffffb18fffff9ada00004e7100006526ffffb18fffff9ada00004e71;
    assign coff[941 ] = 256'hffffb18fffff9ada00004e7100006526ffffb18fffff9ada00004e7100006526;
    assign coff[942 ] = 256'h0000100fffff8103ffffeff100007efd0000100fffff8103ffffeff100007efd;
    assign coff[943 ] = 256'hffff8103ffffeff100007efd0000100fffff8103ffffeff100007efd0000100f;
    assign coff[944 ] = 256'h00007e2fffffea81ffff81d10000157f00007e2fffffea81ffff81d10000157f;
    assign coff[945 ] = 256'hffffea81ffff81d10000157f00007e2fffffea81ffff81d10000157f00007e2f;
    assign coff[946 ] = 256'h00004a06ffff9793ffffb5fa0000686d00004a06ffff9793ffffb5fa0000686d;
    assign coff[947 ] = 256'hffff9793ffffb5fa0000686d00004a06ffff9793ffffb5fa0000686d00004a06;
    assign coff[948 ] = 256'h00006c5affffbbdaffff93a60000442600006c5affffbbdaffff93a600004426;
    assign coff[949 ] = 256'hffffbbdaffff93a60000442600006c5affffbbdaffff93a60000442600006c5a;
    assign coff[950 ] = 256'h00001c6effff8332ffffe39200007cce00001c6effff8332ffffe39200007cce;
    assign coff[951 ] = 256'hffff8332ffffe39200007cce00001c6effff8332ffffe39200007cce00001c6e;
    assign coff[952 ] = 256'h00007790ffffd24dffff887000002db300007790ffffd24dffff887000002db3;
    assign coff[953 ] = 256'hffffd24dffff887000002db300007790ffffd24dffff887000002db300007790;
    assign coff[954 ] = 256'h0000343bffff8b24ffffcbc5000074dc0000343bffff8b24ffffcbc5000074dc;
    assign coff[955 ] = 256'hffff8b24ffffcbc5000074dc0000343bffff8b24ffffcbc5000074dc0000343b;
    assign coff[956 ] = 256'h00005cf9ffffa806ffffa307000057fa00005cf9ffffa806ffffa307000057fa;
    assign coff[957 ] = 256'hffffa806ffffa307000057fa00005cf9ffffa806ffffa307000057fa00005cf9;
    assign coff[958 ] = 256'h00000389ffff800cfffffc7700007ff400000389ffff800cfffffc7700007ff4;
    assign coff[959 ] = 256'hffff800cfffffc7700007ff400000389ffff800cfffffc7700007ff400000389;
    assign coff[960 ] = 256'h00007fddfffffa1dffff8023000005e300007fddfffffa1dffff8023000005e3;
    assign coff[961 ] = 256'hfffffa1dffff8023000005e300007fddfffffa1dffff8023000005e300007fdd;
    assign coff[962 ] = 256'h00005640ffffa16cffffa9c000005e9400005640ffffa16cffffa9c000005e94;
    assign coff[963 ] = 256'hffffa16cffffa9c000005e9400005640ffffa16cffffa9c000005e9400005640;
    assign coff[964 ] = 256'h000073e1ffffc9a1ffff8c1f0000365f000073e1ffffc9a1ffff8c1f0000365f;
    assign coff[965 ] = 256'hffffc9a1ffff8c1f0000365f000073e1ffffc9a1ffff8c1f0000365f000073e1;
    assign coff[966 ] = 256'h00002b7effff879dffffd4820000786300002b7effff879dffffd48200007863;
    assign coff[967 ] = 256'hffff879dffffd4820000786300002b7effff879dffffd4820000786300002b7e;
    assign coff[968 ] = 256'h00007c42ffffe148ffff83be00001eb800007c42ffffe148ffff83be00001eb8;
    assign coff[969 ] = 256'hffffe148ffff83be00001eb800007c42ffffe148ffff83be00001eb800007c42;
    assign coff[970 ] = 256'h00004224ffff926affffbddc00006d9600004224ffff926affffbddc00006d96;
    assign coff[971 ] = 256'hffff926affffbddc00006d9600004224ffff926affffbddc00006d9600004224;
    assign coff[972 ] = 256'h0000670bffffb411ffff98f500004bef0000670bffffb411ffff98f500004bef;
    assign coff[973 ] = 256'hffffb411ffff98f500004bef0000670bffffb411ffff98f500004bef0000670b;
    assign coff[974 ] = 256'h0000132bffff8172ffffecd500007e8e0000132bffff8172ffffecd500007e8e;
    assign coff[975 ] = 256'hffff8172ffffecd500007e8e0000132bffff8172ffffecd500007e8e0000132b;
    assign coff[976 ] = 256'h00007eacffffed9bffff81540000126500007eacffffed9bffff815400001265;
    assign coff[977 ] = 256'hffffed9bffff81540000126500007eacffffed9bffff81540000126500007eac;
    assign coff[978 ] = 256'h00004c91ffff996dffffb36f0000669300004c91ffff996dffffb36f00006693;
    assign coff[979 ] = 256'hffff996dffffb36f0000669300004c91ffff996dffffb36f0000669300004c91;
    assign coff[980 ] = 256'h00006dfeffffbe88ffff92020000417800006dfeffffbe88ffff920200004178;
    assign coff[981 ] = 256'hffffbe88ffff92020000417800006dfeffffbe88ffff92020000417800006dfe;
    assign coff[982 ] = 256'h00001f7bffff83efffffe08500007c1100001f7bffff83efffffe08500007c11;
    assign coff[983 ] = 256'hffff83efffffe08500007c1100001f7bffff83efffffe08500007c1100001f7b;
    assign coff[984 ] = 256'h000078a6ffffd53fffff875a00002ac1000078a6ffffd53fffff875a00002ac1;
    assign coff[985 ] = 256'hffffd53fffff875a00002ac1000078a6ffffd53fffff875a00002ac1000078a6;
    assign coff[986 ] = 256'h00003715ffff8c75ffffc8eb0000738b00003715ffff8c75ffffc8eb0000738b;
    assign coff[987 ] = 256'hffff8c75ffffc8eb0000738b00003715ffff8c75ffffc8eb0000738b00003715;
    assign coff[988 ] = 256'h00005f1bffffaa55ffffa0e5000055ab00005f1bffffaa55ffffa0e5000055ab;
    assign coff[989 ] = 256'hffffaa55ffffa0e5000055ab00005f1bffffaa55ffffa0e5000055ab00005f1b;
    assign coff[990 ] = 256'h000006acffff802dfffff95400007fd3000006acffff802dfffff95400007fd3;
    assign coff[991 ] = 256'hffff802dfffff95400007fd3000006acffff802dfffff95400007fd3000006ac;
    assign coff[992 ] = 256'h00007f6cfffff3d8ffff809400000c2800007f6cfffff3d8ffff809400000c28;
    assign coff[993 ] = 256'hfffff3d8ffff809400000c2800007f6cfffff3d8ffff809400000c2800007f6c;
    assign coff[994 ] = 256'h00005181ffff9d4effffae7f000062b200005181ffff9d4effffae7f000062b2;
    assign coff[995 ] = 256'hffff9d4effffae7f000062b200005181ffff9d4effffae7f000062b200005181;
    assign coff[996 ] = 256'h00007112ffffc402ffff8eee00003bfe00007112ffffc402ffff8eee00003bfe;
    assign coff[997 ] = 256'hffffc402ffff8eee00003bfe00007112ffffc402ffff8eee00003bfe00007112;
    assign coff[998 ] = 256'h00002588ffff85a0ffffda7800007a6000002588ffff85a0ffffda7800007a60;
    assign coff[999 ] = 256'hffff85a0ffffda7800007a6000002588ffff85a0ffffda7800007a6000002588;
    assign coff[1000] = 256'h00007a9affffdb38ffff8566000024c800007a9affffdb38ffff8566000024c8;
    assign coff[1001] = 256'hffffdb38ffff8566000024c800007a9affffdb38ffff8566000024c800007a9a;
    assign coff[1002] = 256'h00003cafffff8f4dffffc351000070b300003cafffff8f4dffffc351000070b3;
    assign coff[1003] = 256'hffff8f4dffffc351000070b300003cafffff8f4dffffc351000070b300003caf;
    assign coff[1004] = 256'h00006332ffffaf1affff9cce000050e600006332ffffaf1affff9cce000050e6;
    assign coff[1005] = 256'hffffaf1affff9cce000050e600006332ffffaf1affff9cce000050e600006332;
    assign coff[1006] = 256'h00000cf0ffff80a8fffff31000007f5800000cf0ffff80a8fffff31000007f58;
    assign coff[1007] = 256'hffff80a8fffff31000007f5800000cf0ffff80a8fffff31000007f5800000cf0;
    assign coff[1008] = 256'h00007d9effffe76affff82620000189600007d9effffe76affff826200001896;
    assign coff[1009] = 256'hffffe76affff82620000189600007d9effffe76affff82620000189600007d9e;
    assign coff[1010] = 256'h00004770ffff95caffffb89000006a3600004770ffff95caffffb89000006a36;
    assign coff[1011] = 256'hffff95caffffb89000006a3600004770ffff95caffffb89000006a3600004770;
    assign coff[1012] = 256'h00006aa5ffffb937ffff955b000046c900006aa5ffffb937ffff955b000046c9;
    assign coff[1013] = 256'hffffb937ffff955b000046c900006aa5ffffb937ffff955b000046c900006aa5;
    assign coff[1014] = 256'h0000195bffff8289ffffe6a500007d770000195bffff8289ffffe6a500007d77;
    assign coff[1015] = 256'hffff8289ffffe6a500007d770000195bffff8289ffffe6a500007d770000195b;
    assign coff[1016] = 256'h00007668ffffcf61ffff89980000309f00007668ffffcf61ffff89980000309f;
    assign coff[1017] = 256'hffffcf61ffff89980000309f00007668ffffcf61ffff89980000309f00007668;
    assign coff[1018] = 256'h00003159ffff89e5ffffcea70000761b00003159ffff89e5ffffcea70000761b;
    assign coff[1019] = 256'hffff89e5ffffcea70000761b00003159ffff89e5ffffcea70000761b00003159;
    assign coff[1020] = 256'h00005ac9ffffa5c5ffffa53700005a3b00005ac9ffffa5c5ffffa53700005a3b;
    assign coff[1021] = 256'hffffa5c5ffffa53700005a3b00005ac9ffffa5c5ffffa53700005a3b00005ac9;
    assign coff[1022] = 256'h00000065ffff8001ffffff9b00007fff00000065ffff8001ffffff9b00007fff;
    assign coff[1023] = 256'hffff8001ffffff9b00007fff00000065ffff8001ffffff9b00007fff00000065;
    assign coff[1024] = 256'h00007fffffffffceffff80010000003200007fffffffffceffff800100000032;
    assign coff[1025] = 256'hffffffceffff80010000003200007fffffffffceffff80010000003200007fff;
    assign coff[1026] = 256'h00005a5fffffa55affffa5a100005aa600005a5fffffa55affffa5a100005aa6;
    assign coff[1027] = 256'hffffa55affffa5a100005aa600005a5fffffa55affffa5a100005aa600005a5f;
    assign coff[1028] = 256'h0000762effffced6ffff89d20000312a0000762effffced6ffff89d20000312a;
    assign coff[1029] = 256'hffffced6ffff89d20000312a0000762effffced6ffff89d20000312a0000762e;
    assign coff[1030] = 256'h000030cdffff89abffffcf3300007655000030cdffff89abffffcf3300007655;
    assign coff[1031] = 256'hffff89abffffcf3300007655000030cdffff89abffffcf3300007655000030cd;
    assign coff[1032] = 256'h00007d81ffffe6d6ffff827f0000192a00007d81ffffe6d6ffff827f0000192a;
    assign coff[1033] = 256'hffffe6d6ffff827f0000192a00007d81ffffe6d6ffff827f0000192a00007d81;
    assign coff[1034] = 256'h000046f3ffff9577ffffb90d00006a89000046f3ffff9577ffffb90d00006a89;
    assign coff[1035] = 256'hffff9577ffffb90d00006a89000046f3ffff9577ffffb90d00006a89000046f3;
    assign coff[1036] = 256'h00006a52ffffb8b9ffff95ae0000474700006a52ffffb8b9ffff95ae00004747;
    assign coff[1037] = 256'hffffb8b9ffff95ae0000474700006a52ffffb8b9ffff95ae0000474700006a52;
    assign coff[1038] = 256'h000018c7ffff826cffffe73900007d94000018c7ffff826cffffe73900007d94;
    assign coff[1039] = 256'hffff826cffffe73900007d94000018c7ffff826cffffe73900007d94000018c7;
    assign coff[1040] = 256'h00007f5dfffff342ffff80a300000cbe00007f5dfffff342ffff80a300000cbe;
    assign coff[1041] = 256'hfffff342ffff80a300000cbe00007f5dfffff342ffff80a300000cbe00007f5d;
    assign coff[1042] = 256'h0000510dffff9ceeffffaef3000063120000510dffff9ceeffffaef300006312;
    assign coff[1043] = 256'hffff9ceeffffaef3000063120000510dffff9ceeffffaef3000063120000510d;
    assign coff[1044] = 256'h000070cbffffc37dffff8f3500003c83000070cbffffc37dffff8f3500003c83;
    assign coff[1045] = 256'hffffc37dffff8f3500003c83000070cbffffc37dffff8f3500003c83000070cb;
    assign coff[1046] = 256'h000024f8ffff8574ffffdb0800007a8c000024f8ffff8574ffffdb0800007a8c;
    assign coff[1047] = 256'hffff8574ffffdb0800007a8c000024f8ffff8574ffffdb0800007a8c000024f8;
    assign coff[1048] = 256'h00007a6effffdaa8ffff85920000255800007a6effffdaa8ffff859200002558;
    assign coff[1049] = 256'hffffdaa8ffff85920000255800007a6effffdaa8ffff85920000255800007a6e;
    assign coff[1050] = 256'h00003c2affff8f06ffffc3d6000070fa00003c2affff8f06ffffc3d6000070fa;
    assign coff[1051] = 256'hffff8f06ffffc3d6000070fa00003c2affff8f06ffffc3d6000070fa00003c2a;
    assign coff[1052] = 256'h000062d2ffffaea5ffff9d2e0000515b000062d2ffffaea5ffff9d2e0000515b;
    assign coff[1053] = 256'hffffaea5ffff9d2e0000515b000062d2ffffaea5ffff9d2e0000515b000062d2;
    assign coff[1054] = 256'h00000c5affff8099fffff3a600007f6700000c5affff8099fffff3a600007f67;
    assign coff[1055] = 256'hffff8099fffff3a600007f6700000c5affff8099fffff3a600007f6700000c5a;
    assign coff[1056] = 256'h00007fd6fffff986ffff802a0000067a00007fd6fffff986ffff802a0000067a;
    assign coff[1057] = 256'hfffff986ffff802a0000067a00007fd6fffff986ffff802a0000067a00007fd6;
    assign coff[1058] = 256'h000055d0ffffa107ffffaa3000005ef9000055d0ffffa107ffffaa3000005ef9;
    assign coff[1059] = 256'hffffa107ffffaa3000005ef9000055d0ffffa107ffffaa3000005ef9000055d0;
    assign coff[1060] = 256'h000073a0ffffc918ffff8c60000036e8000073a0ffffc918ffff8c60000036e8;
    assign coff[1061] = 256'hffffc918ffff8c60000036e8000073a0ffffc918ffff8c60000036e8000073a0;
    assign coff[1062] = 256'h00002af0ffff876bffffd5100000789500002af0ffff876bffffd51000007895;
    assign coff[1063] = 256'hffff876bffffd5100000789500002af0ffff876bffffd5100000789500002af0;
    assign coff[1064] = 256'h00007c1effffe0b5ffff83e200001f4b00007c1effffe0b5ffff83e200001f4b;
    assign coff[1065] = 256'hffffe0b5ffff83e200001f4b00007c1effffe0b5ffff83e200001f4b00007c1e;
    assign coff[1066] = 256'h000041a3ffff921cffffbe5d00006de4000041a3ffff921cffffbe5d00006de4;
    assign coff[1067] = 256'hffff921cffffbe5d00006de4000041a3ffff921cffffbe5d00006de4000041a3;
    assign coff[1068] = 256'h000066b2ffffb398ffff994e00004c68000066b2ffffb398ffff994e00004c68;
    assign coff[1069] = 256'hffffb398ffff994e00004c68000066b2ffffb398ffff994e00004c68000066b2;
    assign coff[1070] = 256'h00001296ffff815bffffed6a00007ea500001296ffff815bffffed6a00007ea5;
    assign coff[1071] = 256'hffff815bffffed6a00007ea500001296ffff815bffffed6a00007ea500001296;
    assign coff[1072] = 256'h00007e96ffffed06ffff816a000012fa00007e96ffffed06ffff816a000012fa;
    assign coff[1073] = 256'hffffed06ffff816a000012fa00007e96ffffed06ffff816a000012fa00007e96;
    assign coff[1074] = 256'h00004c17ffff9913ffffb3e9000066ed00004c17ffff9913ffffb3e9000066ed;
    assign coff[1075] = 256'hffff9913ffffb3e9000066ed00004c17ffff9913ffffb3e9000066ed00004c17;
    assign coff[1076] = 256'h00006db0ffffbe07ffff9250000041f900006db0ffffbe07ffff9250000041f9;
    assign coff[1077] = 256'hffffbe07ffff9250000041f900006db0ffffbe07ffff9250000041f900006db0;
    assign coff[1078] = 256'h00001ee9ffff83caffffe11700007c3600001ee9ffff83caffffe11700007c36;
    assign coff[1079] = 256'hffff83caffffe11700007c3600001ee9ffff83caffffe11700007c3600001ee9;
    assign coff[1080] = 256'h00007874ffffd4b1ffff878c00002b4f00007874ffffd4b1ffff878c00002b4f;
    assign coff[1081] = 256'hffffd4b1ffff878c00002b4f00007874ffffd4b1ffff878c00002b4f00007874;
    assign coff[1082] = 256'h0000368dffff8c35ffffc973000073cb0000368dffff8c35ffffc973000073cb;
    assign coff[1083] = 256'hffff8c35ffffc973000073cb0000368dffff8c35ffffc973000073cb0000368d;
    assign coff[1084] = 256'h00005eb6ffffa9e5ffffa14a0000561b00005eb6ffffa9e5ffffa14a0000561b;
    assign coff[1085] = 256'hffffa9e5ffffa14a0000561b00005eb6ffffa9e5ffffa14a0000561b00005eb6;
    assign coff[1086] = 256'h00000616ffff8025fffff9ea00007fdb00000616ffff8025fffff9ea00007fdb;
    assign coff[1087] = 256'hffff8025fffff9ea00007fdb00000616ffff8025fffff9ea00007fdb00000616;
    assign coff[1088] = 256'h00007ff5fffffcaaffff800b0000035600007ff5fffffcaaffff800b00000356;
    assign coff[1089] = 256'hfffffcaaffff800b0000035600007ff5fffffcaaffff800b0000035600007ff5;
    assign coff[1090] = 256'h0000581effffa329ffffa7e200005cd70000581effffa329ffffa7e200005cd7;
    assign coff[1091] = 256'hffffa329ffffa7e200005cd70000581effffa329ffffa7e200005cd70000581e;
    assign coff[1092] = 256'h000074f0ffffcbf3ffff8b100000340d000074f0ffffcbf3ffff8b100000340d;
    assign coff[1093] = 256'hffffcbf3ffff8b100000340d000074f0ffffcbf3ffff8b100000340d000074f0;
    assign coff[1094] = 256'h00002de2ffff8882ffffd21e0000777e00002de2ffff8882ffffd21e0000777e;
    assign coff[1095] = 256'hffff8882ffffd21e0000777e00002de2ffff8882ffffd21e0000777e00002de2;
    assign coff[1096] = 256'h00007cd9ffffe3c3ffff832700001c3d00007cd9ffffe3c3ffff832700001c3d;
    assign coff[1097] = 256'hffffe3c3ffff832700001c3d00007cd9ffffe3c3ffff832700001c3d00007cd9;
    assign coff[1098] = 256'h00004450ffff93c1ffffbbb000006c3f00004450ffff93c1ffffbbb000006c3f;
    assign coff[1099] = 256'hffff93c1ffffbbb000006c3f00004450ffff93c1ffffbbb000006c3f00004450;
    assign coff[1100] = 256'h0000688affffb623ffff9776000049dd0000688affffb623ffff9776000049dd;
    assign coff[1101] = 256'hffffb623ffff9776000049dd0000688affffb623ffff9776000049dd0000688a;
    assign coff[1102] = 256'h000015b1ffff81daffffea4f00007e26000015b1ffff81daffffea4f00007e26;
    assign coff[1103] = 256'hffff81daffffea4f00007e26000015b1ffff81daffffea4f00007e26000015b1;
    assign coff[1104] = 256'h00007f03fffff023ffff80fd00000fdd00007f03fffff023ffff80fd00000fdd;
    assign coff[1105] = 256'hfffff023ffff80fd00000fdd00007f03fffff023ffff80fd00000fdd00007f03;
    assign coff[1106] = 256'h00004e98ffff9af9ffffb1680000650700004e98ffff9af9ffffb16800006507;
    assign coff[1107] = 256'hffff9af9ffffb1680000650700004e98ffff9af9ffffb1680000650700004e98;
    assign coff[1108] = 256'h00006f46ffffc0bdffff90ba00003f4300006f46ffffc0bdffff90ba00003f43;
    assign coff[1109] = 256'hffffc0bdffff90ba00003f4300006f46ffffc0bdffff90ba00003f4300006f46;
    assign coff[1110] = 256'h000021f3ffff8496ffffde0d00007b6a000021f3ffff8496ffffde0d00007b6a;
    assign coff[1111] = 256'hffff8496ffffde0d00007b6a000021f3ffff8496ffffde0d00007b6a000021f3;
    assign coff[1112] = 256'h0000797affffd7aaffff8686000028560000797affffd7aaffff868600002856;
    assign coff[1113] = 256'hffffd7aaffff8686000028560000797affffd7aaffff8686000028560000797a;
    assign coff[1114] = 256'h00003960ffff8d94ffffc6a00000726c00003960ffff8d94ffffc6a00000726c;
    assign coff[1115] = 256'hffff8d94ffffc6a00000726c00003960ffff8d94ffffc6a00000726c00003960;
    assign coff[1116] = 256'h000060cbffffac3fffff9f35000053c1000060cbffffac3fffff9f35000053c1;
    assign coff[1117] = 256'hffffac3fffff9f35000053c1000060cbffffac3fffff9f35000053c1000060cb;
    assign coff[1118] = 256'h00000938ffff8055fffff6c800007fab00000938ffff8055fffff6c800007fab;
    assign coff[1119] = 256'hffff8055fffff6c800007fab00000938ffff8055fffff6c800007fab00000938;
    assign coff[1120] = 256'h00007fa3fffff663ffff805d0000099d00007fa3fffff663ffff805d0000099d;
    assign coff[1121] = 256'hfffff663ffff805d0000099d00007fa3fffff663ffff805d0000099d00007fa3;
    assign coff[1122] = 256'h00005375ffff9ef3ffffac8b0000610d00005375ffff9ef3ffffac8b0000610d;
    assign coff[1123] = 256'hffff9ef3ffffac8b0000610d00005375ffff9ef3ffffac8b0000610d00005375;
    assign coff[1124] = 256'h0000723fffffc646ffff8dc1000039ba0000723fffffc646ffff8dc1000039ba;
    assign coff[1125] = 256'hffffc646ffff8dc1000039ba0000723fffffc646ffff8dc1000039ba0000723f;
    assign coff[1126] = 256'h000027f7ffff8666ffffd8090000799a000027f7ffff8666ffffd8090000799a;
    assign coff[1127] = 256'hffff8666ffffd8090000799a000027f7ffff8666ffffd8090000799a000027f7;
    assign coff[1128] = 256'h00007b50ffffddacffff84b00000225400007b50ffffddacffff84b000002254;
    assign coff[1129] = 256'hffffddacffff84b00000225400007b50ffffddacffff84b00000225400007b50;
    assign coff[1130] = 256'h00003eecffff9088ffffc11400006f7800003eecffff9088ffffc11400006f78;
    assign coff[1131] = 256'hffff9088ffffc11400006f7800003eecffff9088ffffc11400006f7800003eec;
    assign coff[1132] = 256'h000064caffffb118ffff9b3600004ee8000064caffffb118ffff9b3600004ee8;
    assign coff[1133] = 256'hffffb118ffff9b3600004ee8000064caffffb118ffff9b3600004ee8000064ca;
    assign coff[1134] = 256'h00000f79ffff80f0fffff08700007f1000000f79ffff80f0fffff08700007f10;
    assign coff[1135] = 256'hffff80f0fffff08700007f1000000f79ffff80f0fffff08700007f1000000f79;
    assign coff[1136] = 256'h00007e15ffffe9ecffff81eb0000161400007e15ffffe9ecffff81eb00001614;
    assign coff[1137] = 256'hffffe9ecffff81eb0000161400007e15ffffe9ecffff81eb0000161400007e15;
    assign coff[1138] = 256'h0000498bffff973cffffb675000068c40000498bffff973cffffb675000068c4;
    assign coff[1139] = 256'hffff973cffffb675000068c40000498bffff973cffffb675000068c40000498b;
    assign coff[1140] = 256'h00006c09ffffbb5bffff93f7000044a500006c09ffffbb5bffff93f7000044a5;
    assign coff[1141] = 256'hffffbb5bffff93f7000044a500006c09ffffbb5bffff93f7000044a500006c09;
    assign coff[1142] = 256'h00001bdaffff8311ffffe42600007cef00001bdaffff8311ffffe42600007cef;
    assign coff[1143] = 256'hffff8311ffffe42600007cef00001bdaffff8311ffffe42600007cef00001bda;
    assign coff[1144] = 256'h0000775affffd1c0ffff88a600002e400000775affffd1c0ffff88a600002e40;
    assign coff[1145] = 256'hffffd1c0ffff88a600002e400000775affffd1c0ffff88a600002e400000775a;
    assign coff[1146] = 256'h000033b1ffff8ae7ffffcc4f00007519000033b1ffff8ae7ffffcc4f00007519;
    assign coff[1147] = 256'hffff8ae7ffffcc4f00007519000033b1ffff8ae7ffffcc4f00007519000033b1;
    assign coff[1148] = 256'h00005c91ffffa799ffffa36f0000586700005c91ffffa799ffffa36f00005867;
    assign coff[1149] = 256'hffffa799ffffa36f0000586700005c91ffffa799ffffa36f0000586700005c91;
    assign coff[1150] = 256'h000002f2ffff8009fffffd0e00007ff7000002f2ffff8009fffffd0e00007ff7;
    assign coff[1151] = 256'hffff8009fffffd0e00007ff7000002f2ffff8009fffffd0e00007ff7000002f2;
    assign coff[1152] = 256'h00007ffdfffffe3cffff8003000001c400007ffdfffffe3cffff8003000001c4;
    assign coff[1153] = 256'hfffffe3cffff8003000001c400007ffdfffffe3cffff8003000001c400007ffd;
    assign coff[1154] = 256'h00005940ffffa440ffffa6c000005bc000005940ffffa440ffffa6c000005bc0;
    assign coff[1155] = 256'hffffa440ffffa6c000005bc000005940ffffa440ffffa6c000005bc000005940;
    assign coff[1156] = 256'h00007592ffffcd63ffff8a6e0000329d00007592ffffcd63ffff8a6e0000329d;
    assign coff[1157] = 256'hffffcd63ffff8a6e0000329d00007592ffffcd63ffff8a6e0000329d00007592;
    assign coff[1158] = 256'h00002f59ffff8914ffffd0a7000076ec00002f59ffff8914ffffd0a7000076ec;
    assign coff[1159] = 256'hffff8914ffffd0a7000076ec00002f59ffff8914ffffd0a7000076ec00002f59;
    assign coff[1160] = 256'h00007d2fffffe54cffff82d100001ab400007d2fffffe54cffff82d100001ab4;
    assign coff[1161] = 256'hffffe54cffff82d100001ab400007d2fffffe54cffff82d100001ab400007d2f;
    assign coff[1162] = 256'h000045a3ffff949affffba5d00006b66000045a3ffff949affffba5d00006b66;
    assign coff[1163] = 256'hffff949affffba5d00006b66000045a3ffff949affffba5d00006b66000045a3;
    assign coff[1164] = 256'h00006970ffffb76dffff96900000489300006970ffffb76dffff969000004893;
    assign coff[1165] = 256'hffffb76dffff96900000489300006970ffffb76dffff96900000489300006970;
    assign coff[1166] = 256'h0000173cffff8220ffffe8c400007de00000173cffff8220ffffe8c400007de0;
    assign coff[1167] = 256'hffff8220ffffe8c400007de00000173cffff8220ffffe8c400007de00000173c;
    assign coff[1168] = 256'h00007f33fffff1b2ffff80cd00000e4e00007f33fffff1b2ffff80cd00000e4e;
    assign coff[1169] = 256'hfffff1b2ffff80cd00000e4e00007f33fffff1b2ffff80cd00000e4e00007f33;
    assign coff[1170] = 256'h00004fd4ffff9bf1ffffb02c0000640f00004fd4ffff9bf1ffffb02c0000640f;
    assign coff[1171] = 256'hffff9bf1ffffb02c0000640f00004fd4ffff9bf1ffffb02c0000640f00004fd4;
    assign coff[1172] = 256'h0000700bffffc21cffff8ff500003de40000700bffffc21cffff8ff500003de4;
    assign coff[1173] = 256'hffffc21cffff8ff500003de40000700bffffc21cffff8ff500003de40000700b;
    assign coff[1174] = 256'h00002376ffff8503ffffdc8a00007afd00002376ffff8503ffffdc8a00007afd;
    assign coff[1175] = 256'hffff8503ffffdc8a00007afd00002376ffff8503ffffdc8a00007afd00002376;
    assign coff[1176] = 256'h000079f7ffffd928ffff8609000026d8000079f7ffffd928ffff8609000026d8;
    assign coff[1177] = 256'hffffd928ffff8609000026d8000079f7ffffd928ffff8609000026d8000079f7;
    assign coff[1178] = 256'h00003ac6ffff8e4bffffc53a000071b500003ac6ffff8e4bffffc53a000071b5;
    assign coff[1179] = 256'hffff8e4bffffc53a000071b500003ac6ffff8e4bffffc53a000071b500003ac6;
    assign coff[1180] = 256'h000061d1ffffad70ffff9e2f00005290000061d1ffffad70ffff9e2f00005290;
    assign coff[1181] = 256'hffffad70ffff9e2f00005290000061d1ffffad70ffff9e2f00005290000061d1;
    assign coff[1182] = 256'h00000ac9ffff8075fffff53700007f8b00000ac9ffff8075fffff53700007f8b;
    assign coff[1183] = 256'hffff8075fffff53700007f8b00000ac9ffff8075fffff53700007f8b00000ac9;
    assign coff[1184] = 256'h00007fbffffff7f4ffff80410000080c00007fbffffff7f4ffff80410000080c;
    assign coff[1185] = 256'hfffff7f4ffff80410000080c00007fbffffff7f4ffff80410000080c00007fbf;
    assign coff[1186] = 256'h000054a4ffff9ffbffffab5c00006005000054a4ffff9ffbffffab5c00006005;
    assign coff[1187] = 256'hffff9ffbffffab5c00006005000054a4ffff9ffbffffab5c00006005000054a4;
    assign coff[1188] = 256'h000072f2ffffc7aeffff8d0e00003852000072f2ffffc7aeffff8d0e00003852;
    assign coff[1189] = 256'hffffc7aeffff8d0e00003852000072f2ffffc7aeffff8d0e00003852000072f2;
    assign coff[1190] = 256'h00002974ffff86e6ffffd68c0000791a00002974ffff86e6ffffd68c0000791a;
    assign coff[1191] = 256'hffff86e6ffffd68c0000791a00002974ffff86e6ffffd68c0000791a00002974;
    assign coff[1192] = 256'h00007bb9ffffdf30ffff8447000020d000007bb9ffffdf30ffff8447000020d0;
    assign coff[1193] = 256'hffffdf30ffff8447000020d000007bb9ffffdf30ffff8447000020d000007bb9;
    assign coff[1194] = 256'h00004048ffff9150ffffbfb800006eb000004048ffff9150ffffbfb800006eb0;
    assign coff[1195] = 256'hffff9150ffffbfb800006eb000004048ffff9150ffffbfb800006eb000004048;
    assign coff[1196] = 256'h000065c0ffffb257ffff9a4000004da9000065c0ffffb257ffff9a4000004da9;
    assign coff[1197] = 256'hffffb257ffff9a4000004da9000065c0ffffb257ffff9a4000004da9000065c0;
    assign coff[1198] = 256'h00001108ffff8123ffffeef800007edd00001108ffff8123ffffeef800007edd;
    assign coff[1199] = 256'hffff8123ffffeef800007edd00001108ffff8123ffffeef800007edd00001108;
    assign coff[1200] = 256'h00007e58ffffeb79ffff81a80000148700007e58ffffeb79ffff81a800001487;
    assign coff[1201] = 256'hffffeb79ffff81a80000148700007e58ffffeb79ffff81a80000148700007e58;
    assign coff[1202] = 256'h00004ad3ffff9826ffffb52d000067da00004ad3ffff9826ffffb52d000067da;
    assign coff[1203] = 256'hffff9826ffffb52d000067da00004ad3ffff9826ffffb52d000067da00004ad3;
    assign coff[1204] = 256'h00006cdfffffbcafffff93210000435100006cdfffffbcafffff932100004351;
    assign coff[1205] = 256'hffffbcafffff93210000435100006cdfffffbcafffff93210000435100006cdf;
    assign coff[1206] = 256'h00001d62ffff836bffffe29e00007c9500001d62ffff836bffffe29e00007c95;
    assign coff[1207] = 256'hffff836bffffe29e00007c9500001d62ffff836bffffe29e00007c9500001d62;
    assign coff[1208] = 256'h000077e9ffffd338ffff881700002cc8000077e9ffffd338ffff881700002cc8;
    assign coff[1209] = 256'hffffd338ffff881700002cc8000077e9ffffd338ffff881700002cc8000077e9;
    assign coff[1210] = 256'h00003520ffff8b8bffffcae00000747500003520ffff8b8bffffcae000007475;
    assign coff[1211] = 256'hffff8b8bffffcae00000747500003520ffff8b8bffffcae00000747500003520;
    assign coff[1212] = 256'h00005da5ffffa8bdffffa25b0000574300005da5ffffa8bdffffa25b00005743;
    assign coff[1213] = 256'hffffa8bdffffa25b0000574300005da5ffffa8bdffffa25b0000574300005da5;
    assign coff[1214] = 256'h00000484ffff8014fffffb7c00007fec00000484ffff8014fffffb7c00007fec;
    assign coff[1215] = 256'hffff8014fffffb7c00007fec00000484ffff8014fffffb7c00007fec00000484;
    assign coff[1216] = 256'h00007fe8fffffb18ffff8018000004e800007fe8fffffb18ffff8018000004e8;
    assign coff[1217] = 256'hfffffb18ffff8018000004e800007fe8fffffb18ffff8018000004e800007fe8;
    assign coff[1218] = 256'h000056f9ffffa216ffffa90700005dea000056f9ffffa216ffffa90700005dea;
    assign coff[1219] = 256'hffffa216ffffa90700005dea000056f9ffffa216ffffa90700005dea000056f9;
    assign coff[1220] = 256'h0000744bffffca85ffff8bb50000357b0000744bffffca85ffff8bb50000357b;
    assign coff[1221] = 256'hffffca85ffff8bb50000357b0000744bffffca85ffff8bb50000357b0000744b;
    assign coff[1222] = 256'h00002c6affff87f4ffffd3960000780c00002c6affff87f4ffffd3960000780c;
    assign coff[1223] = 256'hffff87f4ffffd3960000780c00002c6affff87f4ffffd3960000780c00002c6a;
    assign coff[1224] = 256'h00007c7effffe23cffff838200001dc400007c7effffe23cffff838200001dc4;
    assign coff[1225] = 256'hffffe23cffff838200001dc400007c7effffe23cffff838200001dc400007c7e;
    assign coff[1226] = 256'h000042fbffff92ecffffbd0500006d14000042fbffff92ecffffbd0500006d14;
    assign coff[1227] = 256'hffff92ecffffbd0500006d14000042fbffff92ecffffbd0500006d14000042fb;
    assign coff[1228] = 256'h000067a0ffffb4dcffff986000004b24000067a0ffffb4dcffff986000004b24;
    assign coff[1229] = 256'hffffb4dcffff986000004b24000067a0ffffb4dcffff986000004b24000067a0;
    assign coff[1230] = 256'h00001424ffff8198ffffebdc00007e6800001424ffff8198ffffebdc00007e68;
    assign coff[1231] = 256'hffff8198ffffebdc00007e6800001424ffff8198ffffebdc00007e6800001424;
    assign coff[1232] = 256'h00007ecfffffee94ffff81310000116c00007ecfffffee94ffff81310000116c;
    assign coff[1233] = 256'hffffee94ffff81310000116c00007ecfffffee94ffff81310000116c00007ecf;
    assign coff[1234] = 256'h00004d59ffff9a04ffffb2a7000065fc00004d59ffff9a04ffffb2a7000065fc;
    assign coff[1235] = 256'hffff9a04ffffb2a7000065fc00004d59ffff9a04ffffb2a7000065fc00004d59;
    assign coff[1236] = 256'h00006e7dffffbf61ffff91830000409f00006e7dffffbf61ffff91830000409f;
    assign coff[1237] = 256'hffffbf61ffff91830000409f00006e7dffffbf61ffff91830000409f00006e7d;
    assign coff[1238] = 256'h0000206fffff842dffffdf9100007bd30000206fffff842dffffdf9100007bd3;
    assign coff[1239] = 256'hffff842dffffdf9100007bd30000206fffff842dffffdf9100007bd30000206f;
    assign coff[1240] = 256'h000078f9ffffd62dffff8707000029d3000078f9ffffd62dffff8707000029d3;
    assign coff[1241] = 256'hffffd62dffff8707000029d3000078f9ffffd62dffff8707000029d3000078f9;
    assign coff[1242] = 256'h000037f7ffff8ce2ffffc8090000731e000037f7ffff8ce2ffffc8090000731e;
    assign coff[1243] = 256'hffff8ce2ffffc8090000731e000037f7ffff8ce2ffffc8090000731e000037f7;
    assign coff[1244] = 256'h00005fc2ffffab10ffffa03e000054f000005fc2ffffab10ffffa03e000054f0;
    assign coff[1245] = 256'hffffab10ffffa03e000054f000005fc2ffffab10ffffa03e000054f000005fc2;
    assign coff[1246] = 256'h000007a7ffff803bfffff85900007fc5000007a7ffff803bfffff85900007fc5;
    assign coff[1247] = 256'hffff803bfffff85900007fc5000007a7ffff803bfffff85900007fc5000007a7;
    assign coff[1248] = 256'h00007f83fffff4d3ffff807d00000b2d00007f83fffff4d3ffff807d00000b2d;
    assign coff[1249] = 256'hfffff4d3ffff807d00000b2d00007f83fffff4d3ffff807d00000b2d00007f83;
    assign coff[1250] = 256'h00005243ffff9defffffadbd0000621100005243ffff9defffffadbd00006211;
    assign coff[1251] = 256'hffff9defffffadbd0000621100005243ffff9defffffadbd0000621100005243;
    assign coff[1252] = 256'h00007187ffffc4e0ffff8e7900003b2000007187ffffc4e0ffff8e7900003b20;
    assign coff[1253] = 256'hffffc4e0ffff8e7900003b2000007187ffffc4e0ffff8e7900003b2000007187;
    assign coff[1254] = 256'h00002678ffff85ebffffd98800007a1500002678ffff85ebffffd98800007a15;
    assign coff[1255] = 256'hffff85ebffffd98800007a1500002678ffff85ebffffd98800007a1500002678;
    assign coff[1256] = 256'h00007ae1ffffdc29ffff851f000023d700007ae1ffffdc29ffff851f000023d7;
    assign coff[1257] = 256'hffffdc29ffff851f000023d700007ae1ffffdc29ffff851f000023d700007ae1;
    assign coff[1258] = 256'h00003d8cffff8fc5ffffc2740000703b00003d8cffff8fc5ffffc2740000703b;
    assign coff[1259] = 256'hffff8fc5ffffc2740000703b00003d8cffff8fc5ffffc2740000703b00003d8c;
    assign coff[1260] = 256'h000063d0ffffafddffff9c3000005023000063d0ffffafddffff9c3000005023;
    assign coff[1261] = 256'hffffafddffff9c3000005023000063d0ffffafddffff9c3000005023000063d0;
    assign coff[1262] = 256'h00000deaffff80c2fffff21600007f3e00000deaffff80c2fffff21600007f3e;
    assign coff[1263] = 256'hffff80c2fffff21600007f3e00000deaffff80c2fffff21600007f3e00000dea;
    assign coff[1264] = 256'h00007dcdffffe861ffff82330000179f00007dcdffffe861ffff82330000179f;
    assign coff[1265] = 256'hffffe861ffff82330000179f00007dcdffffe861ffff82330000179f00007dcd;
    assign coff[1266] = 256'h00004840ffff9657ffffb7c0000069a900004840ffff9657ffffb7c0000069a9;
    assign coff[1267] = 256'hffff9657ffffb7c0000069a900004840ffff9657ffffb7c0000069a900004840;
    assign coff[1268] = 256'h00006b30ffffba09ffff94d0000045f700006b30ffffba09ffff94d0000045f7;
    assign coff[1269] = 256'hffffba09ffff94d0000045f700006b30ffffba09ffff94d0000045f700006b30;
    assign coff[1270] = 256'h00001a51ffff82bcffffe5af00007d4400001a51ffff82bcffffe5af00007d44;
    assign coff[1271] = 256'hffff82bcffffe5af00007d4400001a51ffff82bcffffe5af00007d4400001a51;
    assign coff[1272] = 256'h000076c7ffffd04affff893900002fb6000076c7ffffd04affff893900002fb6;
    assign coff[1273] = 256'hffffd04affff893900002fb6000076c7ffffd04affff893900002fb6000076c7;
    assign coff[1274] = 256'h00003240ffff8a47ffffcdc0000075b900003240ffff8a47ffffcdc0000075b9;
    assign coff[1275] = 256'hffff8a47ffffcdc0000075b900003240ffff8a47ffffcdc0000075b900003240;
    assign coff[1276] = 256'h00005b7affffa678ffffa4860000598800005b7affffa678ffffa48600005988;
    assign coff[1277] = 256'hffffa678ffffa4860000598800005b7affffa678ffffa4860000598800005b7a;
    assign coff[1278] = 256'h00000160ffff8002fffffea000007ffe00000160ffff8002fffffea000007ffe;
    assign coff[1279] = 256'hffff8002fffffea000007ffe00000160ffff8002fffffea000007ffe00000160;
    assign coff[1280] = 256'h00007fffffffff05ffff8001000000fb00007fffffffff05ffff8001000000fb;
    assign coff[1281] = 256'hffffff05ffff8001000000fb00007fffffffff05ffff8001000000fb00007fff;
    assign coff[1282] = 256'h000059d0ffffa4ccffffa63000005b34000059d0ffffa4ccffffa63000005b34;
    assign coff[1283] = 256'hffffa4ccffffa63000005b34000059d0ffffa4ccffffa63000005b34000059d0;
    assign coff[1284] = 256'h000075e1ffffce1cffff8a1f000031e4000075e1ffffce1cffff8a1f000031e4;
    assign coff[1285] = 256'hffffce1cffff8a1f000031e4000075e1ffffce1cffff8a1f000031e4000075e1;
    assign coff[1286] = 256'h00003013ffff895fffffcfed000076a100003013ffff895fffffcfed000076a1;
    assign coff[1287] = 256'hffff895fffffcfed000076a100003013ffff895fffffcfed000076a100003013;
    assign coff[1288] = 256'h00007d58ffffe611ffff82a8000019ef00007d58ffffe611ffff82a8000019ef;
    assign coff[1289] = 256'hffffe611ffff82a8000019ef00007d58ffffe611ffff82a8000019ef00007d58;
    assign coff[1290] = 256'h0000464bffff9508ffffb9b500006af80000464bffff9508ffffb9b500006af8;
    assign coff[1291] = 256'hffff9508ffffb9b500006af80000464bffff9508ffffb9b500006af80000464b;
    assign coff[1292] = 256'h000069e1ffffb813ffff961f000047ed000069e1ffffb813ffff961f000047ed;
    assign coff[1293] = 256'hffffb813ffff961f000047ed000069e1ffffb813ffff961f000047ed000069e1;
    assign coff[1294] = 256'h00001802ffff8246ffffe7fe00007dba00001802ffff8246ffffe7fe00007dba;
    assign coff[1295] = 256'hffff8246ffffe7fe00007dba00001802ffff8246ffffe7fe00007dba00001802;
    assign coff[1296] = 256'h00007f49fffff27affff80b700000d8600007f49fffff27affff80b700000d86;
    assign coff[1297] = 256'hfffff27affff80b700000d8600007f49fffff27affff80b700000d8600007f49;
    assign coff[1298] = 256'h00005071ffff9c6fffffaf8f0000639100005071ffff9c6fffffaf8f00006391;
    assign coff[1299] = 256'hffff9c6fffffaf8f0000639100005071ffff9c6fffffaf8f0000639100005071;
    assign coff[1300] = 256'h0000706bffffc2ccffff8f9500003d340000706bffffc2ccffff8f9500003d34;
    assign coff[1301] = 256'hffffc2ccffff8f9500003d340000706bffffc2ccffff8f9500003d340000706b;
    assign coff[1302] = 256'h00002437ffff853bffffdbc900007ac500002437ffff853bffffdbc900007ac5;
    assign coff[1303] = 256'hffff853bffffdbc900007ac500002437ffff853bffffdbc900007ac500002437;
    assign coff[1304] = 256'h00007a33ffffd9e8ffff85cd0000261800007a33ffffd9e8ffff85cd00002618;
    assign coff[1305] = 256'hffffd9e8ffff85cd0000261800007a33ffffd9e8ffff85cd0000261800007a33;
    assign coff[1306] = 256'h00003b79ffff8ea8ffffc4870000715800003b79ffff8ea8ffffc48700007158;
    assign coff[1307] = 256'hffff8ea8ffffc4870000715800003b79ffff8ea8ffffc4870000715800003b79;
    assign coff[1308] = 256'h00006252ffffae0bffff9dae000051f500006252ffffae0bffff9dae000051f5;
    assign coff[1309] = 256'hffffae0bffff9dae000051f500006252ffffae0bffff9dae000051f500006252;
    assign coff[1310] = 256'h00000b92ffff8086fffff46e00007f7a00000b92ffff8086fffff46e00007f7a;
    assign coff[1311] = 256'hffff8086fffff46e00007f7a00000b92ffff8086fffff46e00007f7a00000b92;
    assign coff[1312] = 256'h00007fcbfffff8bdffff80350000074300007fcbfffff8bdffff803500000743;
    assign coff[1313] = 256'hfffff8bdffff80350000074300007fcbfffff8bdffff80350000074300007fcb;
    assign coff[1314] = 256'h0000553bffffa080ffffaac500005f800000553bffffa080ffffaac500005f80;
    assign coff[1315] = 256'hffffa080ffffaac500005f800000553bffffa080ffffaac500005f800000553b;
    assign coff[1316] = 256'h0000734affffc863ffff8cb60000379d0000734affffc863ffff8cb60000379d;
    assign coff[1317] = 256'hffffc863ffff8cb60000379d0000734affffc863ffff8cb60000379d0000734a;
    assign coff[1318] = 256'h00002a32ffff8728ffffd5ce000078d800002a32ffff8728ffffd5ce000078d8;
    assign coff[1319] = 256'hffff8728ffffd5ce000078d800002a32ffff8728ffffd5ce000078d800002a32;
    assign coff[1320] = 256'h00007becffffdff2ffff84140000200e00007becffffdff2ffff84140000200e;
    assign coff[1321] = 256'hffffdff2ffff84140000200e00007becffffdff2ffff84140000200e00007bec;
    assign coff[1322] = 256'h000040f6ffff91b6ffffbf0a00006e4a000040f6ffff91b6ffffbf0a00006e4a;
    assign coff[1323] = 256'hffff91b6ffffbf0a00006e4a000040f6ffff91b6ffffbf0a00006e4a000040f6;
    assign coff[1324] = 256'h00006639ffffb2f7ffff99c700004d0900006639ffffb2f7ffff99c700004d09;
    assign coff[1325] = 256'hffffb2f7ffff99c700004d0900006639ffffb2f7ffff99c700004d0900006639;
    assign coff[1326] = 256'h000011cfffff813fffffee3100007ec1000011cfffff813fffffee3100007ec1;
    assign coff[1327] = 256'hffff813fffffee3100007ec1000011cfffff813fffffee3100007ec1000011cf;
    assign coff[1328] = 256'h00007e78ffffec3fffff8188000013c100007e78ffffec3fffff8188000013c1;
    assign coff[1329] = 256'hffffec3fffff8188000013c100007e78ffffec3fffff8188000013c100007e78;
    assign coff[1330] = 256'h00004b75ffff989cffffb48b0000676400004b75ffff989cffffb48b00006764;
    assign coff[1331] = 256'hffff989cffffb48b0000676400004b75ffff989cffffb48b0000676400004b75;
    assign coff[1332] = 256'h00006d48ffffbd5bffff92b8000042a500006d48ffffbd5bffff92b8000042a5;
    assign coff[1333] = 256'hffffbd5bffff92b8000042a500006d48ffffbd5bffff92b8000042a500006d48;
    assign coff[1334] = 256'h00001e26ffff839affffe1da00007c6600001e26ffff839affffe1da00007c66;
    assign coff[1335] = 256'hffff839affffe1da00007c6600001e26ffff839affffe1da00007c6600001e26;
    assign coff[1336] = 256'h0000782fffffd3f4ffff87d100002c0c0000782fffffd3f4ffff87d100002c0c;
    assign coff[1337] = 256'hffffd3f4ffff87d100002c0c0000782fffffd3f4ffff87d100002c0c0000782f;
    assign coff[1338] = 256'h000035d7ffff8bdfffffca2900007421000035d7ffff8bdfffffca2900007421;
    assign coff[1339] = 256'hffff8bdfffffca2900007421000035d7ffff8bdfffffca2900007421000035d7;
    assign coff[1340] = 256'h00005e2effffa951ffffa1d2000056af00005e2effffa951ffffa1d2000056af;
    assign coff[1341] = 256'hffffa951ffffa1d2000056af00005e2effffa951ffffa1d2000056af00005e2e;
    assign coff[1342] = 256'h0000054dffff801cfffffab300007fe40000054dffff801cfffffab300007fe4;
    assign coff[1343] = 256'hffff801cfffffab300007fe40000054dffff801cfffffab300007fe40000054d;
    assign coff[1344] = 256'h00007feffffffbe1ffff80110000041f00007feffffffbe1ffff80110000041f;
    assign coff[1345] = 256'hfffffbe1ffff80110000041f00007feffffffbe1ffff80110000041f00007fef;
    assign coff[1346] = 256'h0000578cffffa29fffffa87400005d610000578cffffa29fffffa87400005d61;
    assign coff[1347] = 256'hffffa29fffffa87400005d610000578cffffa29fffffa87400005d610000578c;
    assign coff[1348] = 256'h0000749effffcb3cffff8b62000034c40000749effffcb3cffff8b62000034c4;
    assign coff[1349] = 256'hffffcb3cffff8b62000034c40000749effffcb3cffff8b62000034c40000749e;
    assign coff[1350] = 256'h00002d26ffff883affffd2da000077c600002d26ffff883affffd2da000077c6;
    assign coff[1351] = 256'hffff883affffd2da000077c600002d26ffff883affffd2da000077c600002d26;
    assign coff[1352] = 256'h00007cacffffe2ffffff835400001d0100007cacffffe2ffffff835400001d01;
    assign coff[1353] = 256'hffffe2ffffff835400001d0100007cacffffe2ffffff835400001d0100007cac;
    assign coff[1354] = 256'h000043a6ffff9356ffffbc5a00006caa000043a6ffff9356ffffbc5a00006caa;
    assign coff[1355] = 256'hffff9356ffffbc5a00006caa000043a6ffff9356ffffbc5a00006caa000043a6;
    assign coff[1356] = 256'h00006815ffffb57fffff97eb00004a8100006815ffffb57fffff97eb00004a81;
    assign coff[1357] = 256'hffffb57fffff97eb00004a8100006815ffffb57fffff97eb00004a8100006815;
    assign coff[1358] = 256'h000014eaffff81b8ffffeb1600007e48000014eaffff81b8ffffeb1600007e48;
    assign coff[1359] = 256'hffff81b8ffffeb1600007e48000014eaffff81b8ffffeb1600007e48000014ea;
    assign coff[1360] = 256'h00007eeaffffef5cffff8116000010a400007eeaffffef5cffff8116000010a4;
    assign coff[1361] = 256'hffffef5cffff8116000010a400007eeaffffef5cffff8116000010a400007eea;
    assign coff[1362] = 256'h00004df9ffff9a7effffb2070000658200004df9ffff9a7effffb20700006582;
    assign coff[1363] = 256'hffff9a7effffb2070000658200004df9ffff9a7effffb2070000658200004df9;
    assign coff[1364] = 256'h00006ee2ffffc00fffff911e00003ff100006ee2ffffc00fffff911e00003ff1;
    assign coff[1365] = 256'hffffc00fffff911e00003ff100006ee2ffffc00fffff911e00003ff100006ee2;
    assign coff[1366] = 256'h00002131ffff8461ffffdecf00007b9f00002131ffff8461ffffdecf00007b9f;
    assign coff[1367] = 256'hffff8461ffffdecf00007b9f00002131ffff8461ffffdecf00007b9f00002131;
    assign coff[1368] = 256'h0000793affffd6ebffff86c6000029150000793affffd6ebffff86c600002915;
    assign coff[1369] = 256'hffffd6ebffff86c6000029150000793affffd6ebffff86c6000029150000793a;
    assign coff[1370] = 256'h000038acffff8d3bffffc754000072c5000038acffff8d3bffffc754000072c5;
    assign coff[1371] = 256'hffff8d3bffffc754000072c5000038acffff8d3bffffc754000072c5000038ac;
    assign coff[1372] = 256'h00006047ffffaba7ffff9fb90000545900006047ffffaba7ffff9fb900005459;
    assign coff[1373] = 256'hffffaba7ffff9fb90000545900006047ffffaba7ffff9fb90000545900006047;
    assign coff[1374] = 256'h00000870ffff8047fffff79000007fb900000870ffff8047fffff79000007fb9;
    assign coff[1375] = 256'hffff8047fffff79000007fb900000870ffff8047fffff79000007fb900000870;
    assign coff[1376] = 256'h00007f94fffff59bffff806c00000a6500007f94fffff59bffff806c00000a65;
    assign coff[1377] = 256'hfffff59bffff806c00000a6500007f94fffff59bffff806c00000a6500007f94;
    assign coff[1378] = 256'h000052dcffff9e70ffffad2400006190000052dcffff9e70ffffad2400006190;
    assign coff[1379] = 256'hffff9e70ffffad2400006190000052dcffff9e70ffffad2400006190000052dc;
    assign coff[1380] = 256'h000071e3ffffc593ffff8e1d00003a6d000071e3ffffc593ffff8e1d00003a6d;
    assign coff[1381] = 256'hffffc593ffff8e1d00003a6d000071e3ffffc593ffff8e1d00003a6d000071e3;
    assign coff[1382] = 256'h00002738ffff8628ffffd8c8000079d800002738ffff8628ffffd8c8000079d8;
    assign coff[1383] = 256'hffff8628ffffd8c8000079d800002738ffff8628ffffd8c8000079d800002738;
    assign coff[1384] = 256'h00007b19ffffdceaffff84e70000231600007b19ffffdceaffff84e700002316;
    assign coff[1385] = 256'hffffdceaffff84e70000231600007b19ffffdceaffff84e70000231600007b19;
    assign coff[1386] = 256'h00003e3cffff9026ffffc1c400006fda00003e3cffff9026ffffc1c400006fda;
    assign coff[1387] = 256'hffff9026ffffc1c400006fda00003e3cffff9026ffffc1c400006fda00003e3c;
    assign coff[1388] = 256'h0000644dffffb07bffff9bb300004f850000644dffffb07bffff9bb300004f85;
    assign coff[1389] = 256'hffffb07bffff9bb300004f850000644dffffb07bffff9bb300004f850000644d;
    assign coff[1390] = 256'h00000eb2ffff80d9fffff14e00007f2700000eb2ffff80d9fffff14e00007f27;
    assign coff[1391] = 256'hffff80d9fffff14e00007f2700000eb2ffff80d9fffff14e00007f2700000eb2;
    assign coff[1392] = 256'h00007df2ffffe926ffff820e000016da00007df2ffffe926ffff820e000016da;
    assign coff[1393] = 256'hffffe926ffff820e000016da00007df2ffffe926ffff820e000016da00007df2;
    assign coff[1394] = 256'h000048e6ffff96c9ffffb71a00006937000048e6ffff96c9ffffb71a00006937;
    assign coff[1395] = 256'hffff96c9ffffb71a00006937000048e6ffff96c9ffffb71a00006937000048e6;
    assign coff[1396] = 256'h00006b9dffffbab1ffff94630000454f00006b9dffffbab1ffff94630000454f;
    assign coff[1397] = 256'hffffbab1ffff94630000454f00006b9dffffbab1ffff94630000454f00006b9d;
    assign coff[1398] = 256'h00001b16ffff82e6ffffe4ea00007d1a00001b16ffff82e6ffffe4ea00007d1a;
    assign coff[1399] = 256'hffff82e6ffffe4ea00007d1a00001b16ffff82e6ffffe4ea00007d1a00001b16;
    assign coff[1400] = 256'h00007711ffffd105ffff88ef00002efb00007711ffffd105ffff88ef00002efb;
    assign coff[1401] = 256'hffffd105ffff88ef00002efb00007711ffffd105ffff88ef00002efb00007711;
    assign coff[1402] = 256'h000032f9ffff8a96ffffcd070000756a000032f9ffff8a96ffffcd070000756a;
    assign coff[1403] = 256'hffff8a96ffffcd070000756a000032f9ffff8a96ffffcd070000756a000032f9;
    assign coff[1404] = 256'h00005c06ffffa708ffffa3fa000058f800005c06ffffa708ffffa3fa000058f8;
    assign coff[1405] = 256'hffffa708ffffa3fa000058f800005c06ffffa708ffffa3fa000058f800005c06;
    assign coff[1406] = 256'h00000229ffff8005fffffdd700007ffb00000229ffff8005fffffdd700007ffb;
    assign coff[1407] = 256'hffff8005fffffdd700007ffb00000229ffff8005fffffdd700007ffb00000229;
    assign coff[1408] = 256'h00007ff9fffffd73ffff80070000028d00007ff9fffffd73ffff80070000028d;
    assign coff[1409] = 256'hfffffd73ffff80070000028d00007ff9fffffd73ffff80070000028d00007ff9;
    assign coff[1410] = 256'h000058b0ffffa3b4ffffa75000005c4c000058b0ffffa3b4ffffa75000005c4c;
    assign coff[1411] = 256'hffffa3b4ffffa75000005c4c000058b0ffffa3b4ffffa75000005c4c000058b0;
    assign coff[1412] = 256'h00007542ffffccabffff8abe0000335500007542ffffccabffff8abe00003355;
    assign coff[1413] = 256'hffffccabffff8abe0000335500007542ffffccabffff8abe0000335500007542;
    assign coff[1414] = 256'h00002e9effff88caffffd1620000773600002e9effff88caffffd16200007736;
    assign coff[1415] = 256'hffff88caffffd1620000773600002e9effff88caffffd1620000773600002e9e;
    assign coff[1416] = 256'h00007d05ffffe488ffff82fb00001b7800007d05ffffe488ffff82fb00001b78;
    assign coff[1417] = 256'hffffe488ffff82fb00001b7800007d05ffffe488ffff82fb00001b7800007d05;
    assign coff[1418] = 256'h000044faffff942dffffbb0600006bd3000044faffff942dffffbb0600006bd3;
    assign coff[1419] = 256'hffff942dffffbb0600006bd3000044faffff942dffffbb0600006bd3000044fa;
    assign coff[1420] = 256'h000068fdffffb6c7ffff970300004939000068fdffffb6c7ffff970300004939;
    assign coff[1421] = 256'hffffb6c7ffff970300004939000068fdffffb6c7ffff970300004939000068fd;
    assign coff[1422] = 256'h00001677ffff81fdffffe98900007e0300001677ffff81fdffffe98900007e03;
    assign coff[1423] = 256'hffff81fdffffe98900007e0300001677ffff81fdffffe98900007e0300001677;
    assign coff[1424] = 256'h00007f1cfffff0ebffff80e400000f1500007f1cfffff0ebffff80e400000f15;
    assign coff[1425] = 256'hfffff0ebffff80e400000f1500007f1cfffff0ebffff80e400000f1500007f1c;
    assign coff[1426] = 256'h00004f37ffff9b75ffffb0c90000648b00004f37ffff9b75ffffb0c90000648b;
    assign coff[1427] = 256'hffff9b75ffffb0c90000648b00004f37ffff9b75ffffb0c90000648b00004f37;
    assign coff[1428] = 256'h00006fa9ffffc16cffff905700003e9400006fa9ffffc16cffff905700003e94;
    assign coff[1429] = 256'hffffc16cffff905700003e9400006fa9ffffc16cffff905700003e9400006fa9;
    assign coff[1430] = 256'h000022b5ffff84ccffffdd4b00007b34000022b5ffff84ccffffdd4b00007b34;
    assign coff[1431] = 256'hffff84ccffffdd4b00007b34000022b5ffff84ccffffdd4b00007b34000022b5;
    assign coff[1432] = 256'h000079b9ffffd869ffff864700002797000079b9ffffd869ffff864700002797;
    assign coff[1433] = 256'hffffd869ffff864700002797000079b9ffffd869ffff864700002797000079b9;
    assign coff[1434] = 256'h00003a13ffff8defffffc5ed0000721100003a13ffff8defffffc5ed00007211;
    assign coff[1435] = 256'hffff8defffffc5ed0000721100003a13ffff8defffffc5ed0000721100003a13;
    assign coff[1436] = 256'h0000614effffacd7ffff9eb2000053290000614effffacd7ffff9eb200005329;
    assign coff[1437] = 256'hffffacd7ffff9eb2000053290000614effffacd7ffff9eb2000053290000614e;
    assign coff[1438] = 256'h00000a01ffff8064fffff5ff00007f9c00000a01ffff8064fffff5ff00007f9c;
    assign coff[1439] = 256'hffff8064fffff5ff00007f9c00000a01ffff8064fffff5ff00007f9c00000a01;
    assign coff[1440] = 256'h00007fb2fffff72cffff804e000008d400007fb2fffff72cffff804e000008d4;
    assign coff[1441] = 256'hfffff72cffff804e000008d400007fb2fffff72cffff804e000008d400007fb2;
    assign coff[1442] = 256'h0000540dffff9f77ffffabf3000060890000540dffff9f77ffffabf300006089;
    assign coff[1443] = 256'hffff9f77ffffabf3000060890000540dffff9f77ffffabf3000060890000540d;
    assign coff[1444] = 256'h00007299ffffc6faffff8d670000390600007299ffffc6faffff8d6700003906;
    assign coff[1445] = 256'hffffc6faffff8d670000390600007299ffffc6faffff8d670000390600007299;
    assign coff[1446] = 256'h000028b6ffff86a5ffffd74a0000795b000028b6ffff86a5ffffd74a0000795b;
    assign coff[1447] = 256'hffff86a5ffffd74a0000795b000028b6ffff86a5ffffd74a0000795b000028b6;
    assign coff[1448] = 256'h00007b85ffffde6effff847b0000219200007b85ffffde6effff847b00002192;
    assign coff[1449] = 256'hffffde6effff847b0000219200007b85ffffde6effff847b0000219200007b85;
    assign coff[1450] = 256'h00003f9affff90ecffffc06600006f1400003f9affff90ecffffc06600006f14;
    assign coff[1451] = 256'hffff90ecffffc06600006f1400003f9affff90ecffffc06600006f1400003f9a;
    assign coff[1452] = 256'h00006545ffffb1b7ffff9abb00004e4900006545ffffb1b7ffff9abb00004e49;
    assign coff[1453] = 256'hffffb1b7ffff9abb00004e4900006545ffffb1b7ffff9abb00004e4900006545;
    assign coff[1454] = 256'h00001041ffff8109ffffefbf00007ef700001041ffff8109ffffefbf00007ef7;
    assign coff[1455] = 256'hffff8109ffffefbf00007ef700001041ffff8109ffffefbf00007ef700001041;
    assign coff[1456] = 256'h00007e37ffffeab3ffff81c90000154d00007e37ffffeab3ffff81c90000154d;
    assign coff[1457] = 256'hffffeab3ffff81c90000154d00007e37ffffeab3ffff81c90000154d00007e37;
    assign coff[1458] = 256'h00004a2fffff97b0ffffb5d10000685000004a2fffff97b0ffffb5d100006850;
    assign coff[1459] = 256'hffff97b0ffffb5d10000685000004a2fffff97b0ffffb5d10000685000004a2f;
    assign coff[1460] = 256'h00006c75ffffbc05ffff938b000043fb00006c75ffffbc05ffff938b000043fb;
    assign coff[1461] = 256'hffffbc05ffff938b000043fb00006c75ffffbc05ffff938b000043fb00006c75;
    assign coff[1462] = 256'h00001c9fffff833effffe36100007cc200001c9fffff833effffe36100007cc2;
    assign coff[1463] = 256'hffff833effffe36100007cc200001c9fffff833effffe36100007cc200001c9f;
    assign coff[1464] = 256'h000077a2ffffd27cffff885e00002d84000077a2ffffd27cffff885e00002d84;
    assign coff[1465] = 256'hffffd27cffff885e00002d84000077a2ffffd27cffff885e00002d84000077a2;
    assign coff[1466] = 256'h00003469ffff8b39ffffcb97000074c700003469ffff8b39ffffcb97000074c7;
    assign coff[1467] = 256'hffff8b39ffffcb97000074c700003469ffff8b39ffffcb97000074c700003469;
    assign coff[1468] = 256'h00005d1cffffa82bffffa2e4000057d500005d1cffffa82bffffa2e4000057d5;
    assign coff[1469] = 256'hffffa82bffffa2e4000057d500005d1cffffa82bffffa2e4000057d500005d1c;
    assign coff[1470] = 256'h000003bbffff800efffffc4500007ff2000003bbffff800efffffc4500007ff2;
    assign coff[1471] = 256'hffff800efffffc4500007ff2000003bbffff800efffffc4500007ff2000003bb;
    assign coff[1472] = 256'h00007fe0fffffa4fffff8020000005b100007fe0fffffa4fffff8020000005b1;
    assign coff[1473] = 256'hfffffa4fffff8020000005b100007fe0fffffa4fffff8020000005b100007fe0;
    assign coff[1474] = 256'h00005665ffffa18effffa99b00005e7200005665ffffa18effffa99b00005e72;
    assign coff[1475] = 256'hffffa18effffa99b00005e7200005665ffffa18effffa99b00005e7200005665;
    assign coff[1476] = 256'h000073f6ffffc9ceffff8c0a00003632000073f6ffffc9ceffff8c0a00003632;
    assign coff[1477] = 256'hffffc9ceffff8c0a00003632000073f6ffffc9ceffff8c0a00003632000073f6;
    assign coff[1478] = 256'h00002badffff87afffffd4530000785100002badffff87afffffd45300007851;
    assign coff[1479] = 256'hffff87afffffd4530000785100002badffff87afffffd4530000785100002bad;
    assign coff[1480] = 256'h00007c4effffe178ffff83b200001e8800007c4effffe178ffff83b200001e88;
    assign coff[1481] = 256'hffffe178ffff83b200001e8800007c4effffe178ffff83b200001e8800007c4e;
    assign coff[1482] = 256'h0000424fffff9284ffffbdb100006d7c0000424fffff9284ffffbdb100006d7c;
    assign coff[1483] = 256'hffff9284ffffbdb100006d7c0000424fffff9284ffffbdb100006d7c0000424f;
    assign coff[1484] = 256'h00006729ffffb439ffff98d700004bc700006729ffffb439ffff98d700004bc7;
    assign coff[1485] = 256'hffffb439ffff98d700004bc700006729ffffb439ffff98d700004bc700006729;
    assign coff[1486] = 256'h0000135dffff8179ffffeca300007e870000135dffff8179ffffeca300007e87;
    assign coff[1487] = 256'hffff8179ffffeca300007e870000135dffff8179ffffeca300007e870000135d;
    assign coff[1488] = 256'h00007eb3ffffedcdffff814d0000123300007eb3ffffedcdffff814d00001233;
    assign coff[1489] = 256'hffffedcdffff814d0000123300007eb3ffffedcdffff814d0000123300007eb3;
    assign coff[1490] = 256'h00004cb9ffff998bffffb3470000667500004cb9ffff998bffffb34700006675;
    assign coff[1491] = 256'hffff998bffffb3470000667500004cb9ffff998bffffb3470000667500004cb9;
    assign coff[1492] = 256'h00006e17ffffbeb3ffff91e90000414d00006e17ffffbeb3ffff91e90000414d;
    assign coff[1493] = 256'hffffbeb3ffff91e90000414d00006e17ffffbeb3ffff91e90000414d00006e17;
    assign coff[1494] = 256'h00001facffff83fbffffe05400007c0500001facffff83fbffffe05400007c05;
    assign coff[1495] = 256'hffff83fbffffe05400007c0500001facffff83fbffffe05400007c0500001fac;
    assign coff[1496] = 256'h000078b7ffffd56fffff874900002a91000078b7ffffd56fffff874900002a91;
    assign coff[1497] = 256'hffffd56fffff874900002a91000078b7ffffd56fffff874900002a91000078b7;
    assign coff[1498] = 256'h00003742ffff8c8bffffc8be0000737500003742ffff8c8bffffc8be00007375;
    assign coff[1499] = 256'hffff8c8bffffc8be0000737500003742ffff8c8bffffc8be0000737500003742;
    assign coff[1500] = 256'h00005f3cffffaa7affffa0c40000558600005f3cffffaa7affffa0c400005586;
    assign coff[1501] = 256'hffffaa7affffa0c40000558600005f3cffffaa7affffa0c40000558600005f3c;
    assign coff[1502] = 256'h000006deffff802ffffff92200007fd1000006deffff802ffffff92200007fd1;
    assign coff[1503] = 256'hffff802ffffff92200007fd1000006deffff802ffffff92200007fd1000006de;
    assign coff[1504] = 256'h00007f71fffff40affff808f00000bf600007f71fffff40affff808f00000bf6;
    assign coff[1505] = 256'hfffff40affff808f00000bf600007f71fffff40affff808f00000bf600007f71;
    assign coff[1506] = 256'h000051a8ffff9d6effffae5800006292000051a8ffff9d6effffae5800006292;
    assign coff[1507] = 256'hffff9d6effffae5800006292000051a8ffff9d6effffae5800006292000051a8;
    assign coff[1508] = 256'h0000712affffc42effff8ed600003bd20000712affffc42effff8ed600003bd2;
    assign coff[1509] = 256'hffffc42effff8ed600003bd20000712affffc42effff8ed600003bd20000712a;
    assign coff[1510] = 256'h000025b8ffff85afffffda4800007a51000025b8ffff85afffffda4800007a51;
    assign coff[1511] = 256'hffff85afffffda4800007a51000025b8ffff85afffffda4800007a51000025b8;
    assign coff[1512] = 256'h00007aa8ffffdb68ffff85580000249800007aa8ffffdb68ffff855800002498;
    assign coff[1513] = 256'hffffdb68ffff85580000249800007aa8ffffdb68ffff85580000249800007aa8;
    assign coff[1514] = 256'h00003cdcffff8f65ffffc3240000709b00003cdcffff8f65ffffc3240000709b;
    assign coff[1515] = 256'hffff8f65ffffc3240000709b00003cdcffff8f65ffffc3240000709b00003cdc;
    assign coff[1516] = 256'h00006351ffffaf41ffff9caf000050bf00006351ffffaf41ffff9caf000050bf;
    assign coff[1517] = 256'hffffaf41ffff9caf000050bf00006351ffffaf41ffff9caf000050bf00006351;
    assign coff[1518] = 256'h00000d22ffff80adfffff2de00007f5300000d22ffff80adfffff2de00007f53;
    assign coff[1519] = 256'hffff80adfffff2de00007f5300000d22ffff80adfffff2de00007f5300000d22;
    assign coff[1520] = 256'h00007da7ffffe79bffff82590000186500007da7ffffe79bffff825900001865;
    assign coff[1521] = 256'hffffe79bffff82590000186500007da7ffffe79bffff82590000186500007da7;
    assign coff[1522] = 256'h0000479affff95e6ffffb86600006a1a0000479affff95e6ffffb86600006a1a;
    assign coff[1523] = 256'hffff95e6ffffb86600006a1a0000479affff95e6ffffb86600006a1a0000479a;
    assign coff[1524] = 256'h00006ac1ffffb961ffff953f0000469f00006ac1ffffb961ffff953f0000469f;
    assign coff[1525] = 256'hffffb961ffff953f0000469f00006ac1ffffb961ffff953f0000469f00006ac1;
    assign coff[1526] = 256'h0000198dffff8293ffffe67300007d6d0000198dffff8293ffffe67300007d6d;
    assign coff[1527] = 256'hffff8293ffffe67300007d6d0000198dffff8293ffffe67300007d6d0000198d;
    assign coff[1528] = 256'h0000767bffffcf90ffff8985000030700000767bffffcf90ffff898500003070;
    assign coff[1529] = 256'hffffcf90ffff8985000030700000767bffffcf90ffff8985000030700000767b;
    assign coff[1530] = 256'h00003187ffff89f8ffffce790000760800003187ffff89f8ffffce7900007608;
    assign coff[1531] = 256'hffff89f8ffffce790000760800003187ffff89f8ffffce790000760800003187;
    assign coff[1532] = 256'h00005aedffffa5e8ffffa51300005a1800005aedffffa5e8ffffa51300005a18;
    assign coff[1533] = 256'hffffa5e8ffffa51300005a1800005aedffffa5e8ffffa51300005a1800005aed;
    assign coff[1534] = 256'h00000097ffff8001ffffff6900007fff00000097ffff8001ffffff6900007fff;
    assign coff[1535] = 256'hffff8001ffffff6900007fff00000097ffff8001ffffff6900007fff00000097;
    assign coff[1536] = 256'h00007fffffffff69ffff80010000009700007fffffffff69ffff800100000097;
    assign coff[1537] = 256'hffffff69ffff80010000009700007fffffffff69ffff80010000009700007fff;
    assign coff[1538] = 256'h00005a18ffffa513ffffa5e800005aed00005a18ffffa513ffffa5e800005aed;
    assign coff[1539] = 256'hffffa513ffffa5e800005aed00005a18ffffa513ffffa5e800005aed00005a18;
    assign coff[1540] = 256'h00007608ffffce79ffff89f80000318700007608ffffce79ffff89f800003187;
    assign coff[1541] = 256'hffffce79ffff89f80000318700007608ffffce79ffff89f80000318700007608;
    assign coff[1542] = 256'h00003070ffff8985ffffcf900000767b00003070ffff8985ffffcf900000767b;
    assign coff[1543] = 256'hffff8985ffffcf900000767b00003070ffff8985ffffcf900000767b00003070;
    assign coff[1544] = 256'h00007d6dffffe673ffff82930000198d00007d6dffffe673ffff82930000198d;
    assign coff[1545] = 256'hffffe673ffff82930000198d00007d6dffffe673ffff82930000198d00007d6d;
    assign coff[1546] = 256'h0000469fffff953fffffb96100006ac10000469fffff953fffffb96100006ac1;
    assign coff[1547] = 256'hffff953fffffb96100006ac10000469fffff953fffffb96100006ac10000469f;
    assign coff[1548] = 256'h00006a1affffb866ffff95e60000479a00006a1affffb866ffff95e60000479a;
    assign coff[1549] = 256'hffffb866ffff95e60000479a00006a1affffb866ffff95e60000479a00006a1a;
    assign coff[1550] = 256'h00001865ffff8259ffffe79b00007da700001865ffff8259ffffe79b00007da7;
    assign coff[1551] = 256'hffff8259ffffe79b00007da700001865ffff8259ffffe79b00007da700001865;
    assign coff[1552] = 256'h00007f53fffff2deffff80ad00000d2200007f53fffff2deffff80ad00000d22;
    assign coff[1553] = 256'hfffff2deffff80ad00000d2200007f53fffff2deffff80ad00000d2200007f53;
    assign coff[1554] = 256'h000050bfffff9cafffffaf4100006351000050bfffff9cafffffaf4100006351;
    assign coff[1555] = 256'hffff9cafffffaf4100006351000050bfffff9cafffffaf4100006351000050bf;
    assign coff[1556] = 256'h0000709bffffc324ffff8f6500003cdc0000709bffffc324ffff8f6500003cdc;
    assign coff[1557] = 256'hffffc324ffff8f6500003cdc0000709bffffc324ffff8f6500003cdc0000709b;
    assign coff[1558] = 256'h00002498ffff8558ffffdb6800007aa800002498ffff8558ffffdb6800007aa8;
    assign coff[1559] = 256'hffff8558ffffdb6800007aa800002498ffff8558ffffdb6800007aa800002498;
    assign coff[1560] = 256'h00007a51ffffda48ffff85af000025b800007a51ffffda48ffff85af000025b8;
    assign coff[1561] = 256'hffffda48ffff85af000025b800007a51ffffda48ffff85af000025b800007a51;
    assign coff[1562] = 256'h00003bd2ffff8ed6ffffc42e0000712a00003bd2ffff8ed6ffffc42e0000712a;
    assign coff[1563] = 256'hffff8ed6ffffc42e0000712a00003bd2ffff8ed6ffffc42e0000712a00003bd2;
    assign coff[1564] = 256'h00006292ffffae58ffff9d6e000051a800006292ffffae58ffff9d6e000051a8;
    assign coff[1565] = 256'hffffae58ffff9d6e000051a800006292ffffae58ffff9d6e000051a800006292;
    assign coff[1566] = 256'h00000bf6ffff808ffffff40a00007f7100000bf6ffff808ffffff40a00007f71;
    assign coff[1567] = 256'hffff808ffffff40a00007f7100000bf6ffff808ffffff40a00007f7100000bf6;
    assign coff[1568] = 256'h00007fd1fffff922ffff802f000006de00007fd1fffff922ffff802f000006de;
    assign coff[1569] = 256'hfffff922ffff802f000006de00007fd1fffff922ffff802f000006de00007fd1;
    assign coff[1570] = 256'h00005586ffffa0c4ffffaa7a00005f3c00005586ffffa0c4ffffaa7a00005f3c;
    assign coff[1571] = 256'hffffa0c4ffffaa7a00005f3c00005586ffffa0c4ffffaa7a00005f3c00005586;
    assign coff[1572] = 256'h00007375ffffc8beffff8c8b0000374200007375ffffc8beffff8c8b00003742;
    assign coff[1573] = 256'hffffc8beffff8c8b0000374200007375ffffc8beffff8c8b0000374200007375;
    assign coff[1574] = 256'h00002a91ffff8749ffffd56f000078b700002a91ffff8749ffffd56f000078b7;
    assign coff[1575] = 256'hffff8749ffffd56f000078b700002a91ffff8749ffffd56f000078b700002a91;
    assign coff[1576] = 256'h00007c05ffffe054ffff83fb00001fac00007c05ffffe054ffff83fb00001fac;
    assign coff[1577] = 256'hffffe054ffff83fb00001fac00007c05ffffe054ffff83fb00001fac00007c05;
    assign coff[1578] = 256'h0000414dffff91e9ffffbeb300006e170000414dffff91e9ffffbeb300006e17;
    assign coff[1579] = 256'hffff91e9ffffbeb300006e170000414dffff91e9ffffbeb300006e170000414d;
    assign coff[1580] = 256'h00006675ffffb347ffff998b00004cb900006675ffffb347ffff998b00004cb9;
    assign coff[1581] = 256'hffffb347ffff998b00004cb900006675ffffb347ffff998b00004cb900006675;
    assign coff[1582] = 256'h00001233ffff814dffffedcd00007eb300001233ffff814dffffedcd00007eb3;
    assign coff[1583] = 256'hffff814dffffedcd00007eb300001233ffff814dffffedcd00007eb300001233;
    assign coff[1584] = 256'h00007e87ffffeca3ffff81790000135d00007e87ffffeca3ffff81790000135d;
    assign coff[1585] = 256'hffffeca3ffff81790000135d00007e87ffffeca3ffff81790000135d00007e87;
    assign coff[1586] = 256'h00004bc7ffff98d7ffffb4390000672900004bc7ffff98d7ffffb43900006729;
    assign coff[1587] = 256'hffff98d7ffffb4390000672900004bc7ffff98d7ffffb4390000672900004bc7;
    assign coff[1588] = 256'h00006d7cffffbdb1ffff92840000424f00006d7cffffbdb1ffff92840000424f;
    assign coff[1589] = 256'hffffbdb1ffff92840000424f00006d7cffffbdb1ffff92840000424f00006d7c;
    assign coff[1590] = 256'h00001e88ffff83b2ffffe17800007c4e00001e88ffff83b2ffffe17800007c4e;
    assign coff[1591] = 256'hffff83b2ffffe17800007c4e00001e88ffff83b2ffffe17800007c4e00001e88;
    assign coff[1592] = 256'h00007851ffffd453ffff87af00002bad00007851ffffd453ffff87af00002bad;
    assign coff[1593] = 256'hffffd453ffff87af00002bad00007851ffffd453ffff87af00002bad00007851;
    assign coff[1594] = 256'h00003632ffff8c0affffc9ce000073f600003632ffff8c0affffc9ce000073f6;
    assign coff[1595] = 256'hffff8c0affffc9ce000073f600003632ffff8c0affffc9ce000073f600003632;
    assign coff[1596] = 256'h00005e72ffffa99bffffa18e0000566500005e72ffffa99bffffa18e00005665;
    assign coff[1597] = 256'hffffa99bffffa18e0000566500005e72ffffa99bffffa18e0000566500005e72;
    assign coff[1598] = 256'h000005b1ffff8020fffffa4f00007fe0000005b1ffff8020fffffa4f00007fe0;
    assign coff[1599] = 256'hffff8020fffffa4f00007fe0000005b1ffff8020fffffa4f00007fe0000005b1;
    assign coff[1600] = 256'h00007ff2fffffc45ffff800e000003bb00007ff2fffffc45ffff800e000003bb;
    assign coff[1601] = 256'hfffffc45ffff800e000003bb00007ff2fffffc45ffff800e000003bb00007ff2;
    assign coff[1602] = 256'h000057d5ffffa2e4ffffa82b00005d1c000057d5ffffa2e4ffffa82b00005d1c;
    assign coff[1603] = 256'hffffa2e4ffffa82b00005d1c000057d5ffffa2e4ffffa82b00005d1c000057d5;
    assign coff[1604] = 256'h000074c7ffffcb97ffff8b3900003469000074c7ffffcb97ffff8b3900003469;
    assign coff[1605] = 256'hffffcb97ffff8b3900003469000074c7ffffcb97ffff8b3900003469000074c7;
    assign coff[1606] = 256'h00002d84ffff885effffd27c000077a200002d84ffff885effffd27c000077a2;
    assign coff[1607] = 256'hffff885effffd27c000077a200002d84ffff885effffd27c000077a200002d84;
    assign coff[1608] = 256'h00007cc2ffffe361ffff833e00001c9f00007cc2ffffe361ffff833e00001c9f;
    assign coff[1609] = 256'hffffe361ffff833e00001c9f00007cc2ffffe361ffff833e00001c9f00007cc2;
    assign coff[1610] = 256'h000043fbffff938bffffbc0500006c75000043fbffff938bffffbc0500006c75;
    assign coff[1611] = 256'hffff938bffffbc0500006c75000043fbffff938bffffbc0500006c75000043fb;
    assign coff[1612] = 256'h00006850ffffb5d1ffff97b000004a2f00006850ffffb5d1ffff97b000004a2f;
    assign coff[1613] = 256'hffffb5d1ffff97b000004a2f00006850ffffb5d1ffff97b000004a2f00006850;
    assign coff[1614] = 256'h0000154dffff81c9ffffeab300007e370000154dffff81c9ffffeab300007e37;
    assign coff[1615] = 256'hffff81c9ffffeab300007e370000154dffff81c9ffffeab300007e370000154d;
    assign coff[1616] = 256'h00007ef7ffffefbfffff81090000104100007ef7ffffefbfffff810900001041;
    assign coff[1617] = 256'hffffefbfffff81090000104100007ef7ffffefbfffff81090000104100007ef7;
    assign coff[1618] = 256'h00004e49ffff9abbffffb1b70000654500004e49ffff9abbffffb1b700006545;
    assign coff[1619] = 256'hffff9abbffffb1b70000654500004e49ffff9abbffffb1b70000654500004e49;
    assign coff[1620] = 256'h00006f14ffffc066ffff90ec00003f9a00006f14ffffc066ffff90ec00003f9a;
    assign coff[1621] = 256'hffffc066ffff90ec00003f9a00006f14ffffc066ffff90ec00003f9a00006f14;
    assign coff[1622] = 256'h00002192ffff847bffffde6e00007b8500002192ffff847bffffde6e00007b85;
    assign coff[1623] = 256'hffff847bffffde6e00007b8500002192ffff847bffffde6e00007b8500002192;
    assign coff[1624] = 256'h0000795bffffd74affff86a5000028b60000795bffffd74affff86a5000028b6;
    assign coff[1625] = 256'hffffd74affff86a5000028b60000795bffffd74affff86a5000028b60000795b;
    assign coff[1626] = 256'h00003906ffff8d67ffffc6fa0000729900003906ffff8d67ffffc6fa00007299;
    assign coff[1627] = 256'hffff8d67ffffc6fa0000729900003906ffff8d67ffffc6fa0000729900003906;
    assign coff[1628] = 256'h00006089ffffabf3ffff9f770000540d00006089ffffabf3ffff9f770000540d;
    assign coff[1629] = 256'hffffabf3ffff9f770000540d00006089ffffabf3ffff9f770000540d00006089;
    assign coff[1630] = 256'h000008d4ffff804efffff72c00007fb2000008d4ffff804efffff72c00007fb2;
    assign coff[1631] = 256'hffff804efffff72c00007fb2000008d4ffff804efffff72c00007fb2000008d4;
    assign coff[1632] = 256'h00007f9cfffff5ffffff806400000a0100007f9cfffff5ffffff806400000a01;
    assign coff[1633] = 256'hfffff5ffffff806400000a0100007f9cfffff5ffffff806400000a0100007f9c;
    assign coff[1634] = 256'h00005329ffff9eb2ffffacd70000614e00005329ffff9eb2ffffacd70000614e;
    assign coff[1635] = 256'hffff9eb2ffffacd70000614e00005329ffff9eb2ffffacd70000614e00005329;
    assign coff[1636] = 256'h00007211ffffc5edffff8def00003a1300007211ffffc5edffff8def00003a13;
    assign coff[1637] = 256'hffffc5edffff8def00003a1300007211ffffc5edffff8def00003a1300007211;
    assign coff[1638] = 256'h00002797ffff8647ffffd869000079b900002797ffff8647ffffd869000079b9;
    assign coff[1639] = 256'hffff8647ffffd869000079b900002797ffff8647ffffd869000079b900002797;
    assign coff[1640] = 256'h00007b34ffffdd4bffff84cc000022b500007b34ffffdd4bffff84cc000022b5;
    assign coff[1641] = 256'hffffdd4bffff84cc000022b500007b34ffffdd4bffff84cc000022b500007b34;
    assign coff[1642] = 256'h00003e94ffff9057ffffc16c00006fa900003e94ffff9057ffffc16c00006fa9;
    assign coff[1643] = 256'hffff9057ffffc16c00006fa900003e94ffff9057ffffc16c00006fa900003e94;
    assign coff[1644] = 256'h0000648bffffb0c9ffff9b7500004f370000648bffffb0c9ffff9b7500004f37;
    assign coff[1645] = 256'hffffb0c9ffff9b7500004f370000648bffffb0c9ffff9b7500004f370000648b;
    assign coff[1646] = 256'h00000f15ffff80e4fffff0eb00007f1c00000f15ffff80e4fffff0eb00007f1c;
    assign coff[1647] = 256'hffff80e4fffff0eb00007f1c00000f15ffff80e4fffff0eb00007f1c00000f15;
    assign coff[1648] = 256'h00007e03ffffe989ffff81fd0000167700007e03ffffe989ffff81fd00001677;
    assign coff[1649] = 256'hffffe989ffff81fd0000167700007e03ffffe989ffff81fd0000167700007e03;
    assign coff[1650] = 256'h00004939ffff9703ffffb6c7000068fd00004939ffff9703ffffb6c7000068fd;
    assign coff[1651] = 256'hffff9703ffffb6c7000068fd00004939ffff9703ffffb6c7000068fd00004939;
    assign coff[1652] = 256'h00006bd3ffffbb06ffff942d000044fa00006bd3ffffbb06ffff942d000044fa;
    assign coff[1653] = 256'hffffbb06ffff942d000044fa00006bd3ffffbb06ffff942d000044fa00006bd3;
    assign coff[1654] = 256'h00001b78ffff82fbffffe48800007d0500001b78ffff82fbffffe48800007d05;
    assign coff[1655] = 256'hffff82fbffffe48800007d0500001b78ffff82fbffffe48800007d0500001b78;
    assign coff[1656] = 256'h00007736ffffd162ffff88ca00002e9e00007736ffffd162ffff88ca00002e9e;
    assign coff[1657] = 256'hffffd162ffff88ca00002e9e00007736ffffd162ffff88ca00002e9e00007736;
    assign coff[1658] = 256'h00003355ffff8abeffffccab0000754200003355ffff8abeffffccab00007542;
    assign coff[1659] = 256'hffff8abeffffccab0000754200003355ffff8abeffffccab0000754200003355;
    assign coff[1660] = 256'h00005c4cffffa750ffffa3b4000058b000005c4cffffa750ffffa3b4000058b0;
    assign coff[1661] = 256'hffffa750ffffa3b4000058b000005c4cffffa750ffffa3b4000058b000005c4c;
    assign coff[1662] = 256'h0000028dffff8007fffffd7300007ff90000028dffff8007fffffd7300007ff9;
    assign coff[1663] = 256'hffff8007fffffd7300007ff90000028dffff8007fffffd7300007ff90000028d;
    assign coff[1664] = 256'h00007ffbfffffdd7ffff80050000022900007ffbfffffdd7ffff800500000229;
    assign coff[1665] = 256'hfffffdd7ffff80050000022900007ffbfffffdd7ffff80050000022900007ffb;
    assign coff[1666] = 256'h000058f8ffffa3faffffa70800005c06000058f8ffffa3faffffa70800005c06;
    assign coff[1667] = 256'hffffa3faffffa70800005c06000058f8ffffa3faffffa70800005c06000058f8;
    assign coff[1668] = 256'h0000756affffcd07ffff8a96000032f90000756affffcd07ffff8a96000032f9;
    assign coff[1669] = 256'hffffcd07ffff8a96000032f90000756affffcd07ffff8a96000032f90000756a;
    assign coff[1670] = 256'h00002efbffff88efffffd1050000771100002efbffff88efffffd10500007711;
    assign coff[1671] = 256'hffff88efffffd1050000771100002efbffff88efffffd1050000771100002efb;
    assign coff[1672] = 256'h00007d1affffe4eaffff82e600001b1600007d1affffe4eaffff82e600001b16;
    assign coff[1673] = 256'hffffe4eaffff82e600001b1600007d1affffe4eaffff82e600001b1600007d1a;
    assign coff[1674] = 256'h0000454fffff9463ffffbab100006b9d0000454fffff9463ffffbab100006b9d;
    assign coff[1675] = 256'hffff9463ffffbab100006b9d0000454fffff9463ffffbab100006b9d0000454f;
    assign coff[1676] = 256'h00006937ffffb71affff96c9000048e600006937ffffb71affff96c9000048e6;
    assign coff[1677] = 256'hffffb71affff96c9000048e600006937ffffb71affff96c9000048e600006937;
    assign coff[1678] = 256'h000016daffff820effffe92600007df2000016daffff820effffe92600007df2;
    assign coff[1679] = 256'hffff820effffe92600007df2000016daffff820effffe92600007df2000016da;
    assign coff[1680] = 256'h00007f27fffff14effff80d900000eb200007f27fffff14effff80d900000eb2;
    assign coff[1681] = 256'hfffff14effff80d900000eb200007f27fffff14effff80d900000eb200007f27;
    assign coff[1682] = 256'h00004f85ffff9bb3ffffb07b0000644d00004f85ffff9bb3ffffb07b0000644d;
    assign coff[1683] = 256'hffff9bb3ffffb07b0000644d00004f85ffff9bb3ffffb07b0000644d00004f85;
    assign coff[1684] = 256'h00006fdaffffc1c4ffff902600003e3c00006fdaffffc1c4ffff902600003e3c;
    assign coff[1685] = 256'hffffc1c4ffff902600003e3c00006fdaffffc1c4ffff902600003e3c00006fda;
    assign coff[1686] = 256'h00002316ffff84e7ffffdcea00007b1900002316ffff84e7ffffdcea00007b19;
    assign coff[1687] = 256'hffff84e7ffffdcea00007b1900002316ffff84e7ffffdcea00007b1900002316;
    assign coff[1688] = 256'h000079d8ffffd8c8ffff862800002738000079d8ffffd8c8ffff862800002738;
    assign coff[1689] = 256'hffffd8c8ffff862800002738000079d8ffffd8c8ffff862800002738000079d8;
    assign coff[1690] = 256'h00003a6dffff8e1dffffc593000071e300003a6dffff8e1dffffc593000071e3;
    assign coff[1691] = 256'hffff8e1dffffc593000071e300003a6dffff8e1dffffc593000071e300003a6d;
    assign coff[1692] = 256'h00006190ffffad24ffff9e70000052dc00006190ffffad24ffff9e70000052dc;
    assign coff[1693] = 256'hffffad24ffff9e70000052dc00006190ffffad24ffff9e70000052dc00006190;
    assign coff[1694] = 256'h00000a65ffff806cfffff59b00007f9400000a65ffff806cfffff59b00007f94;
    assign coff[1695] = 256'hffff806cfffff59b00007f9400000a65ffff806cfffff59b00007f9400000a65;
    assign coff[1696] = 256'h00007fb9fffff790ffff80470000087000007fb9fffff790ffff804700000870;
    assign coff[1697] = 256'hfffff790ffff80470000087000007fb9fffff790ffff80470000087000007fb9;
    assign coff[1698] = 256'h00005459ffff9fb9ffffaba70000604700005459ffff9fb9ffffaba700006047;
    assign coff[1699] = 256'hffff9fb9ffffaba70000604700005459ffff9fb9ffffaba70000604700005459;
    assign coff[1700] = 256'h000072c5ffffc754ffff8d3b000038ac000072c5ffffc754ffff8d3b000038ac;
    assign coff[1701] = 256'hffffc754ffff8d3b000038ac000072c5ffffc754ffff8d3b000038ac000072c5;
    assign coff[1702] = 256'h00002915ffff86c6ffffd6eb0000793a00002915ffff86c6ffffd6eb0000793a;
    assign coff[1703] = 256'hffff86c6ffffd6eb0000793a00002915ffff86c6ffffd6eb0000793a00002915;
    assign coff[1704] = 256'h00007b9fffffdecfffff84610000213100007b9fffffdecfffff846100002131;
    assign coff[1705] = 256'hffffdecfffff84610000213100007b9fffffdecfffff84610000213100007b9f;
    assign coff[1706] = 256'h00003ff1ffff911effffc00f00006ee200003ff1ffff911effffc00f00006ee2;
    assign coff[1707] = 256'hffff911effffc00f00006ee200003ff1ffff911effffc00f00006ee200003ff1;
    assign coff[1708] = 256'h00006582ffffb207ffff9a7e00004df900006582ffffb207ffff9a7e00004df9;
    assign coff[1709] = 256'hffffb207ffff9a7e00004df900006582ffffb207ffff9a7e00004df900006582;
    assign coff[1710] = 256'h000010a4ffff8116ffffef5c00007eea000010a4ffff8116ffffef5c00007eea;
    assign coff[1711] = 256'hffff8116ffffef5c00007eea000010a4ffff8116ffffef5c00007eea000010a4;
    assign coff[1712] = 256'h00007e48ffffeb16ffff81b8000014ea00007e48ffffeb16ffff81b8000014ea;
    assign coff[1713] = 256'hffffeb16ffff81b8000014ea00007e48ffffeb16ffff81b8000014ea00007e48;
    assign coff[1714] = 256'h00004a81ffff97ebffffb57f0000681500004a81ffff97ebffffb57f00006815;
    assign coff[1715] = 256'hffff97ebffffb57f0000681500004a81ffff97ebffffb57f0000681500004a81;
    assign coff[1716] = 256'h00006caaffffbc5affff9356000043a600006caaffffbc5affff9356000043a6;
    assign coff[1717] = 256'hffffbc5affff9356000043a600006caaffffbc5affff9356000043a600006caa;
    assign coff[1718] = 256'h00001d01ffff8354ffffe2ff00007cac00001d01ffff8354ffffe2ff00007cac;
    assign coff[1719] = 256'hffff8354ffffe2ff00007cac00001d01ffff8354ffffe2ff00007cac00001d01;
    assign coff[1720] = 256'h000077c6ffffd2daffff883a00002d26000077c6ffffd2daffff883a00002d26;
    assign coff[1721] = 256'hffffd2daffff883a00002d26000077c6ffffd2daffff883a00002d26000077c6;
    assign coff[1722] = 256'h000034c4ffff8b62ffffcb3c0000749e000034c4ffff8b62ffffcb3c0000749e;
    assign coff[1723] = 256'hffff8b62ffffcb3c0000749e000034c4ffff8b62ffffcb3c0000749e000034c4;
    assign coff[1724] = 256'h00005d61ffffa874ffffa29f0000578c00005d61ffffa874ffffa29f0000578c;
    assign coff[1725] = 256'hffffa874ffffa29f0000578c00005d61ffffa874ffffa29f0000578c00005d61;
    assign coff[1726] = 256'h0000041fffff8011fffffbe100007fef0000041fffff8011fffffbe100007fef;
    assign coff[1727] = 256'hffff8011fffffbe100007fef0000041fffff8011fffffbe100007fef0000041f;
    assign coff[1728] = 256'h00007fe4fffffab3ffff801c0000054d00007fe4fffffab3ffff801c0000054d;
    assign coff[1729] = 256'hfffffab3ffff801c0000054d00007fe4fffffab3ffff801c0000054d00007fe4;
    assign coff[1730] = 256'h000056afffffa1d2ffffa95100005e2e000056afffffa1d2ffffa95100005e2e;
    assign coff[1731] = 256'hffffa1d2ffffa95100005e2e000056afffffa1d2ffffa95100005e2e000056af;
    assign coff[1732] = 256'h00007421ffffca29ffff8bdf000035d700007421ffffca29ffff8bdf000035d7;
    assign coff[1733] = 256'hffffca29ffff8bdf000035d700007421ffffca29ffff8bdf000035d700007421;
    assign coff[1734] = 256'h00002c0cffff87d1ffffd3f40000782f00002c0cffff87d1ffffd3f40000782f;
    assign coff[1735] = 256'hffff87d1ffffd3f40000782f00002c0cffff87d1ffffd3f40000782f00002c0c;
    assign coff[1736] = 256'h00007c66ffffe1daffff839a00001e2600007c66ffffe1daffff839a00001e26;
    assign coff[1737] = 256'hffffe1daffff839a00001e2600007c66ffffe1daffff839a00001e2600007c66;
    assign coff[1738] = 256'h000042a5ffff92b8ffffbd5b00006d48000042a5ffff92b8ffffbd5b00006d48;
    assign coff[1739] = 256'hffff92b8ffffbd5b00006d48000042a5ffff92b8ffffbd5b00006d48000042a5;
    assign coff[1740] = 256'h00006764ffffb48bffff989c00004b7500006764ffffb48bffff989c00004b75;
    assign coff[1741] = 256'hffffb48bffff989c00004b7500006764ffffb48bffff989c00004b7500006764;
    assign coff[1742] = 256'h000013c1ffff8188ffffec3f00007e78000013c1ffff8188ffffec3f00007e78;
    assign coff[1743] = 256'hffff8188ffffec3f00007e78000013c1ffff8188ffffec3f00007e78000013c1;
    assign coff[1744] = 256'h00007ec1ffffee31ffff813f000011cf00007ec1ffffee31ffff813f000011cf;
    assign coff[1745] = 256'hffffee31ffff813f000011cf00007ec1ffffee31ffff813f000011cf00007ec1;
    assign coff[1746] = 256'h00004d09ffff99c7ffffb2f70000663900004d09ffff99c7ffffb2f700006639;
    assign coff[1747] = 256'hffff99c7ffffb2f70000663900004d09ffff99c7ffffb2f70000663900004d09;
    assign coff[1748] = 256'h00006e4affffbf0affff91b6000040f600006e4affffbf0affff91b6000040f6;
    assign coff[1749] = 256'hffffbf0affff91b6000040f600006e4affffbf0affff91b6000040f600006e4a;
    assign coff[1750] = 256'h0000200effff8414ffffdff200007bec0000200effff8414ffffdff200007bec;
    assign coff[1751] = 256'hffff8414ffffdff200007bec0000200effff8414ffffdff200007bec0000200e;
    assign coff[1752] = 256'h000078d8ffffd5ceffff872800002a32000078d8ffffd5ceffff872800002a32;
    assign coff[1753] = 256'hffffd5ceffff872800002a32000078d8ffffd5ceffff872800002a32000078d8;
    assign coff[1754] = 256'h0000379dffff8cb6ffffc8630000734a0000379dffff8cb6ffffc8630000734a;
    assign coff[1755] = 256'hffff8cb6ffffc8630000734a0000379dffff8cb6ffffc8630000734a0000379d;
    assign coff[1756] = 256'h00005f80ffffaac5ffffa0800000553b00005f80ffffaac5ffffa0800000553b;
    assign coff[1757] = 256'hffffaac5ffffa0800000553b00005f80ffffaac5ffffa0800000553b00005f80;
    assign coff[1758] = 256'h00000743ffff8035fffff8bd00007fcb00000743ffff8035fffff8bd00007fcb;
    assign coff[1759] = 256'hffff8035fffff8bd00007fcb00000743ffff8035fffff8bd00007fcb00000743;
    assign coff[1760] = 256'h00007f7afffff46effff808600000b9200007f7afffff46effff808600000b92;
    assign coff[1761] = 256'hfffff46effff808600000b9200007f7afffff46effff808600000b9200007f7a;
    assign coff[1762] = 256'h000051f5ffff9daeffffae0b00006252000051f5ffff9daeffffae0b00006252;
    assign coff[1763] = 256'hffff9daeffffae0b00006252000051f5ffff9daeffffae0b00006252000051f5;
    assign coff[1764] = 256'h00007158ffffc487ffff8ea800003b7900007158ffffc487ffff8ea800003b79;
    assign coff[1765] = 256'hffffc487ffff8ea800003b7900007158ffffc487ffff8ea800003b7900007158;
    assign coff[1766] = 256'h00002618ffff85cdffffd9e800007a3300002618ffff85cdffffd9e800007a33;
    assign coff[1767] = 256'hffff85cdffffd9e800007a3300002618ffff85cdffffd9e800007a3300002618;
    assign coff[1768] = 256'h00007ac5ffffdbc9ffff853b0000243700007ac5ffffdbc9ffff853b00002437;
    assign coff[1769] = 256'hffffdbc9ffff853b0000243700007ac5ffffdbc9ffff853b0000243700007ac5;
    assign coff[1770] = 256'h00003d34ffff8f95ffffc2cc0000706b00003d34ffff8f95ffffc2cc0000706b;
    assign coff[1771] = 256'hffff8f95ffffc2cc0000706b00003d34ffff8f95ffffc2cc0000706b00003d34;
    assign coff[1772] = 256'h00006391ffffaf8fffff9c6f0000507100006391ffffaf8fffff9c6f00005071;
    assign coff[1773] = 256'hffffaf8fffff9c6f0000507100006391ffffaf8fffff9c6f0000507100006391;
    assign coff[1774] = 256'h00000d86ffff80b7fffff27a00007f4900000d86ffff80b7fffff27a00007f49;
    assign coff[1775] = 256'hffff80b7fffff27a00007f4900000d86ffff80b7fffff27a00007f4900000d86;
    assign coff[1776] = 256'h00007dbaffffe7feffff82460000180200007dbaffffe7feffff824600001802;
    assign coff[1777] = 256'hffffe7feffff82460000180200007dbaffffe7feffff82460000180200007dba;
    assign coff[1778] = 256'h000047edffff961fffffb813000069e1000047edffff961fffffb813000069e1;
    assign coff[1779] = 256'hffff961fffffb813000069e1000047edffff961fffffb813000069e1000047ed;
    assign coff[1780] = 256'h00006af8ffffb9b5ffff95080000464b00006af8ffffb9b5ffff95080000464b;
    assign coff[1781] = 256'hffffb9b5ffff95080000464b00006af8ffffb9b5ffff95080000464b00006af8;
    assign coff[1782] = 256'h000019efffff82a8ffffe61100007d58000019efffff82a8ffffe61100007d58;
    assign coff[1783] = 256'hffff82a8ffffe61100007d58000019efffff82a8ffffe61100007d58000019ef;
    assign coff[1784] = 256'h000076a1ffffcfedffff895f00003013000076a1ffffcfedffff895f00003013;
    assign coff[1785] = 256'hffffcfedffff895f00003013000076a1ffffcfedffff895f00003013000076a1;
    assign coff[1786] = 256'h000031e4ffff8a1fffffce1c000075e1000031e4ffff8a1fffffce1c000075e1;
    assign coff[1787] = 256'hffff8a1fffffce1c000075e1000031e4ffff8a1fffffce1c000075e1000031e4;
    assign coff[1788] = 256'h00005b34ffffa630ffffa4cc000059d000005b34ffffa630ffffa4cc000059d0;
    assign coff[1789] = 256'hffffa630ffffa4cc000059d000005b34ffffa630ffffa4cc000059d000005b34;
    assign coff[1790] = 256'h000000fbffff8001ffffff0500007fff000000fbffff8001ffffff0500007fff;
    assign coff[1791] = 256'hffff8001ffffff0500007fff000000fbffff8001ffffff0500007fff000000fb;
    assign coff[1792] = 256'h00007ffefffffea0ffff80020000016000007ffefffffea0ffff800200000160;
    assign coff[1793] = 256'hfffffea0ffff80020000016000007ffefffffea0ffff80020000016000007ffe;
    assign coff[1794] = 256'h00005988ffffa486ffffa67800005b7a00005988ffffa486ffffa67800005b7a;
    assign coff[1795] = 256'hffffa486ffffa67800005b7a00005988ffffa486ffffa67800005b7a00005988;
    assign coff[1796] = 256'h000075b9ffffcdc0ffff8a4700003240000075b9ffffcdc0ffff8a4700003240;
    assign coff[1797] = 256'hffffcdc0ffff8a4700003240000075b9ffffcdc0ffff8a4700003240000075b9;
    assign coff[1798] = 256'h00002fb6ffff8939ffffd04a000076c700002fb6ffff8939ffffd04a000076c7;
    assign coff[1799] = 256'hffff8939ffffd04a000076c700002fb6ffff8939ffffd04a000076c700002fb6;
    assign coff[1800] = 256'h00007d44ffffe5afffff82bc00001a5100007d44ffffe5afffff82bc00001a51;
    assign coff[1801] = 256'hffffe5afffff82bc00001a5100007d44ffffe5afffff82bc00001a5100007d44;
    assign coff[1802] = 256'h000045f7ffff94d0ffffba0900006b30000045f7ffff94d0ffffba0900006b30;
    assign coff[1803] = 256'hffff94d0ffffba0900006b30000045f7ffff94d0ffffba0900006b30000045f7;
    assign coff[1804] = 256'h000069a9ffffb7c0ffff965700004840000069a9ffffb7c0ffff965700004840;
    assign coff[1805] = 256'hffffb7c0ffff965700004840000069a9ffffb7c0ffff965700004840000069a9;
    assign coff[1806] = 256'h0000179fffff8233ffffe86100007dcd0000179fffff8233ffffe86100007dcd;
    assign coff[1807] = 256'hffff8233ffffe86100007dcd0000179fffff8233ffffe86100007dcd0000179f;
    assign coff[1808] = 256'h00007f3efffff216ffff80c200000dea00007f3efffff216ffff80c200000dea;
    assign coff[1809] = 256'hfffff216ffff80c200000dea00007f3efffff216ffff80c200000dea00007f3e;
    assign coff[1810] = 256'h00005023ffff9c30ffffafdd000063d000005023ffff9c30ffffafdd000063d0;
    assign coff[1811] = 256'hffff9c30ffffafdd000063d000005023ffff9c30ffffafdd000063d000005023;
    assign coff[1812] = 256'h0000703bffffc274ffff8fc500003d8c0000703bffffc274ffff8fc500003d8c;
    assign coff[1813] = 256'hffffc274ffff8fc500003d8c0000703bffffc274ffff8fc500003d8c0000703b;
    assign coff[1814] = 256'h000023d7ffff851fffffdc2900007ae1000023d7ffff851fffffdc2900007ae1;
    assign coff[1815] = 256'hffff851fffffdc2900007ae1000023d7ffff851fffffdc2900007ae1000023d7;
    assign coff[1816] = 256'h00007a15ffffd988ffff85eb0000267800007a15ffffd988ffff85eb00002678;
    assign coff[1817] = 256'hffffd988ffff85eb0000267800007a15ffffd988ffff85eb0000267800007a15;
    assign coff[1818] = 256'h00003b20ffff8e79ffffc4e00000718700003b20ffff8e79ffffc4e000007187;
    assign coff[1819] = 256'hffff8e79ffffc4e00000718700003b20ffff8e79ffffc4e00000718700003b20;
    assign coff[1820] = 256'h00006211ffffadbdffff9def0000524300006211ffffadbdffff9def00005243;
    assign coff[1821] = 256'hffffadbdffff9def0000524300006211ffffadbdffff9def0000524300006211;
    assign coff[1822] = 256'h00000b2dffff807dfffff4d300007f8300000b2dffff807dfffff4d300007f83;
    assign coff[1823] = 256'hffff807dfffff4d300007f8300000b2dffff807dfffff4d300007f8300000b2d;
    assign coff[1824] = 256'h00007fc5fffff859ffff803b000007a700007fc5fffff859ffff803b000007a7;
    assign coff[1825] = 256'hfffff859ffff803b000007a700007fc5fffff859ffff803b000007a700007fc5;
    assign coff[1826] = 256'h000054f0ffffa03effffab1000005fc2000054f0ffffa03effffab1000005fc2;
    assign coff[1827] = 256'hffffa03effffab1000005fc2000054f0ffffa03effffab1000005fc2000054f0;
    assign coff[1828] = 256'h0000731effffc809ffff8ce2000037f70000731effffc809ffff8ce2000037f7;
    assign coff[1829] = 256'hffffc809ffff8ce2000037f70000731effffc809ffff8ce2000037f70000731e;
    assign coff[1830] = 256'h000029d3ffff8707ffffd62d000078f9000029d3ffff8707ffffd62d000078f9;
    assign coff[1831] = 256'hffff8707ffffd62d000078f9000029d3ffff8707ffffd62d000078f9000029d3;
    assign coff[1832] = 256'h00007bd3ffffdf91ffff842d0000206f00007bd3ffffdf91ffff842d0000206f;
    assign coff[1833] = 256'hffffdf91ffff842d0000206f00007bd3ffffdf91ffff842d0000206f00007bd3;
    assign coff[1834] = 256'h0000409fffff9183ffffbf6100006e7d0000409fffff9183ffffbf6100006e7d;
    assign coff[1835] = 256'hffff9183ffffbf6100006e7d0000409fffff9183ffffbf6100006e7d0000409f;
    assign coff[1836] = 256'h000065fcffffb2a7ffff9a0400004d59000065fcffffb2a7ffff9a0400004d59;
    assign coff[1837] = 256'hffffb2a7ffff9a0400004d59000065fcffffb2a7ffff9a0400004d59000065fc;
    assign coff[1838] = 256'h0000116cffff8131ffffee9400007ecf0000116cffff8131ffffee9400007ecf;
    assign coff[1839] = 256'hffff8131ffffee9400007ecf0000116cffff8131ffffee9400007ecf0000116c;
    assign coff[1840] = 256'h00007e68ffffebdcffff81980000142400007e68ffffebdcffff819800001424;
    assign coff[1841] = 256'hffffebdcffff81980000142400007e68ffffebdcffff81980000142400007e68;
    assign coff[1842] = 256'h00004b24ffff9860ffffb4dc000067a000004b24ffff9860ffffb4dc000067a0;
    assign coff[1843] = 256'hffff9860ffffb4dc000067a000004b24ffff9860ffffb4dc000067a000004b24;
    assign coff[1844] = 256'h00006d14ffffbd05ffff92ec000042fb00006d14ffffbd05ffff92ec000042fb;
    assign coff[1845] = 256'hffffbd05ffff92ec000042fb00006d14ffffbd05ffff92ec000042fb00006d14;
    assign coff[1846] = 256'h00001dc4ffff8382ffffe23c00007c7e00001dc4ffff8382ffffe23c00007c7e;
    assign coff[1847] = 256'hffff8382ffffe23c00007c7e00001dc4ffff8382ffffe23c00007c7e00001dc4;
    assign coff[1848] = 256'h0000780cffffd396ffff87f400002c6a0000780cffffd396ffff87f400002c6a;
    assign coff[1849] = 256'hffffd396ffff87f400002c6a0000780cffffd396ffff87f400002c6a0000780c;
    assign coff[1850] = 256'h0000357bffff8bb5ffffca850000744b0000357bffff8bb5ffffca850000744b;
    assign coff[1851] = 256'hffff8bb5ffffca850000744b0000357bffff8bb5ffffca850000744b0000357b;
    assign coff[1852] = 256'h00005deaffffa907ffffa216000056f900005deaffffa907ffffa216000056f9;
    assign coff[1853] = 256'hffffa907ffffa216000056f900005deaffffa907ffffa216000056f900005dea;
    assign coff[1854] = 256'h000004e8ffff8018fffffb1800007fe8000004e8ffff8018fffffb1800007fe8;
    assign coff[1855] = 256'hffff8018fffffb1800007fe8000004e8ffff8018fffffb1800007fe8000004e8;
    assign coff[1856] = 256'h00007fecfffffb7cffff80140000048400007fecfffffb7cffff801400000484;
    assign coff[1857] = 256'hfffffb7cffff80140000048400007fecfffffb7cffff80140000048400007fec;
    assign coff[1858] = 256'h00005743ffffa25bffffa8bd00005da500005743ffffa25bffffa8bd00005da5;
    assign coff[1859] = 256'hffffa25bffffa8bd00005da500005743ffffa25bffffa8bd00005da500005743;
    assign coff[1860] = 256'h00007475ffffcae0ffff8b8b0000352000007475ffffcae0ffff8b8b00003520;
    assign coff[1861] = 256'hffffcae0ffff8b8b0000352000007475ffffcae0ffff8b8b0000352000007475;
    assign coff[1862] = 256'h00002cc8ffff8817ffffd338000077e900002cc8ffff8817ffffd338000077e9;
    assign coff[1863] = 256'hffff8817ffffd338000077e900002cc8ffff8817ffffd338000077e900002cc8;
    assign coff[1864] = 256'h00007c95ffffe29effff836b00001d6200007c95ffffe29effff836b00001d62;
    assign coff[1865] = 256'hffffe29effff836b00001d6200007c95ffffe29effff836b00001d6200007c95;
    assign coff[1866] = 256'h00004351ffff9321ffffbcaf00006cdf00004351ffff9321ffffbcaf00006cdf;
    assign coff[1867] = 256'hffff9321ffffbcaf00006cdf00004351ffff9321ffffbcaf00006cdf00004351;
    assign coff[1868] = 256'h000067daffffb52dffff982600004ad3000067daffffb52dffff982600004ad3;
    assign coff[1869] = 256'hffffb52dffff982600004ad3000067daffffb52dffff982600004ad3000067da;
    assign coff[1870] = 256'h00001487ffff81a8ffffeb7900007e5800001487ffff81a8ffffeb7900007e58;
    assign coff[1871] = 256'hffff81a8ffffeb7900007e5800001487ffff81a8ffffeb7900007e5800001487;
    assign coff[1872] = 256'h00007eddffffeef8ffff81230000110800007eddffffeef8ffff812300001108;
    assign coff[1873] = 256'hffffeef8ffff81230000110800007eddffffeef8ffff81230000110800007edd;
    assign coff[1874] = 256'h00004da9ffff9a40ffffb257000065c000004da9ffff9a40ffffb257000065c0;
    assign coff[1875] = 256'hffff9a40ffffb257000065c000004da9ffff9a40ffffb257000065c000004da9;
    assign coff[1876] = 256'h00006eb0ffffbfb8ffff91500000404800006eb0ffffbfb8ffff915000004048;
    assign coff[1877] = 256'hffffbfb8ffff91500000404800006eb0ffffbfb8ffff91500000404800006eb0;
    assign coff[1878] = 256'h000020d0ffff8447ffffdf3000007bb9000020d0ffff8447ffffdf3000007bb9;
    assign coff[1879] = 256'hffff8447ffffdf3000007bb9000020d0ffff8447ffffdf3000007bb9000020d0;
    assign coff[1880] = 256'h0000791affffd68cffff86e6000029740000791affffd68cffff86e600002974;
    assign coff[1881] = 256'hffffd68cffff86e6000029740000791affffd68cffff86e6000029740000791a;
    assign coff[1882] = 256'h00003852ffff8d0effffc7ae000072f200003852ffff8d0effffc7ae000072f2;
    assign coff[1883] = 256'hffff8d0effffc7ae000072f200003852ffff8d0effffc7ae000072f200003852;
    assign coff[1884] = 256'h00006005ffffab5cffff9ffb000054a400006005ffffab5cffff9ffb000054a4;
    assign coff[1885] = 256'hffffab5cffff9ffb000054a400006005ffffab5cffff9ffb000054a400006005;
    assign coff[1886] = 256'h0000080cffff8041fffff7f400007fbf0000080cffff8041fffff7f400007fbf;
    assign coff[1887] = 256'hffff8041fffff7f400007fbf0000080cffff8041fffff7f400007fbf0000080c;
    assign coff[1888] = 256'h00007f8bfffff537ffff807500000ac900007f8bfffff537ffff807500000ac9;
    assign coff[1889] = 256'hfffff537ffff807500000ac900007f8bfffff537ffff807500000ac900007f8b;
    assign coff[1890] = 256'h00005290ffff9e2fffffad70000061d100005290ffff9e2fffffad70000061d1;
    assign coff[1891] = 256'hffff9e2fffffad70000061d100005290ffff9e2fffffad70000061d100005290;
    assign coff[1892] = 256'h000071b5ffffc53affff8e4b00003ac6000071b5ffffc53affff8e4b00003ac6;
    assign coff[1893] = 256'hffffc53affff8e4b00003ac6000071b5ffffc53affff8e4b00003ac6000071b5;
    assign coff[1894] = 256'h000026d8ffff8609ffffd928000079f7000026d8ffff8609ffffd928000079f7;
    assign coff[1895] = 256'hffff8609ffffd928000079f7000026d8ffff8609ffffd928000079f7000026d8;
    assign coff[1896] = 256'h00007afdffffdc8affff85030000237600007afdffffdc8affff850300002376;
    assign coff[1897] = 256'hffffdc8affff85030000237600007afdffffdc8affff85030000237600007afd;
    assign coff[1898] = 256'h00003de4ffff8ff5ffffc21c0000700b00003de4ffff8ff5ffffc21c0000700b;
    assign coff[1899] = 256'hffff8ff5ffffc21c0000700b00003de4ffff8ff5ffffc21c0000700b00003de4;
    assign coff[1900] = 256'h0000640fffffb02cffff9bf100004fd40000640fffffb02cffff9bf100004fd4;
    assign coff[1901] = 256'hffffb02cffff9bf100004fd40000640fffffb02cffff9bf100004fd40000640f;
    assign coff[1902] = 256'h00000e4effff80cdfffff1b200007f3300000e4effff80cdfffff1b200007f33;
    assign coff[1903] = 256'hffff80cdfffff1b200007f3300000e4effff80cdfffff1b200007f3300000e4e;
    assign coff[1904] = 256'h00007de0ffffe8c4ffff82200000173c00007de0ffffe8c4ffff82200000173c;
    assign coff[1905] = 256'hffffe8c4ffff82200000173c00007de0ffffe8c4ffff82200000173c00007de0;
    assign coff[1906] = 256'h00004893ffff9690ffffb76d0000697000004893ffff9690ffffb76d00006970;
    assign coff[1907] = 256'hffff9690ffffb76d0000697000004893ffff9690ffffb76d0000697000004893;
    assign coff[1908] = 256'h00006b66ffffba5dffff949a000045a300006b66ffffba5dffff949a000045a3;
    assign coff[1909] = 256'hffffba5dffff949a000045a300006b66ffffba5dffff949a000045a300006b66;
    assign coff[1910] = 256'h00001ab4ffff82d1ffffe54c00007d2f00001ab4ffff82d1ffffe54c00007d2f;
    assign coff[1911] = 256'hffff82d1ffffe54c00007d2f00001ab4ffff82d1ffffe54c00007d2f00001ab4;
    assign coff[1912] = 256'h000076ecffffd0a7ffff891400002f59000076ecffffd0a7ffff891400002f59;
    assign coff[1913] = 256'hffffd0a7ffff891400002f59000076ecffffd0a7ffff891400002f59000076ec;
    assign coff[1914] = 256'h0000329dffff8a6effffcd63000075920000329dffff8a6effffcd6300007592;
    assign coff[1915] = 256'hffff8a6effffcd63000075920000329dffff8a6effffcd63000075920000329d;
    assign coff[1916] = 256'h00005bc0ffffa6c0ffffa4400000594000005bc0ffffa6c0ffffa44000005940;
    assign coff[1917] = 256'hffffa6c0ffffa4400000594000005bc0ffffa6c0ffffa4400000594000005bc0;
    assign coff[1918] = 256'h000001c4ffff8003fffffe3c00007ffd000001c4ffff8003fffffe3c00007ffd;
    assign coff[1919] = 256'hffff8003fffffe3c00007ffd000001c4ffff8003fffffe3c00007ffd000001c4;
    assign coff[1920] = 256'h00007ff7fffffd0effff8009000002f200007ff7fffffd0effff8009000002f2;
    assign coff[1921] = 256'hfffffd0effff8009000002f200007ff7fffffd0effff8009000002f200007ff7;
    assign coff[1922] = 256'h00005867ffffa36fffffa79900005c9100005867ffffa36fffffa79900005c91;
    assign coff[1923] = 256'hffffa36fffffa79900005c9100005867ffffa36fffffa79900005c9100005867;
    assign coff[1924] = 256'h00007519ffffcc4fffff8ae7000033b100007519ffffcc4fffff8ae7000033b1;
    assign coff[1925] = 256'hffffcc4fffff8ae7000033b100007519ffffcc4fffff8ae7000033b100007519;
    assign coff[1926] = 256'h00002e40ffff88a6ffffd1c00000775a00002e40ffff88a6ffffd1c00000775a;
    assign coff[1927] = 256'hffff88a6ffffd1c00000775a00002e40ffff88a6ffffd1c00000775a00002e40;
    assign coff[1928] = 256'h00007cefffffe426ffff831100001bda00007cefffffe426ffff831100001bda;
    assign coff[1929] = 256'hffffe426ffff831100001bda00007cefffffe426ffff831100001bda00007cef;
    assign coff[1930] = 256'h000044a5ffff93f7ffffbb5b00006c09000044a5ffff93f7ffffbb5b00006c09;
    assign coff[1931] = 256'hffff93f7ffffbb5b00006c09000044a5ffff93f7ffffbb5b00006c09000044a5;
    assign coff[1932] = 256'h000068c4ffffb675ffff973c0000498b000068c4ffffb675ffff973c0000498b;
    assign coff[1933] = 256'hffffb675ffff973c0000498b000068c4ffffb675ffff973c0000498b000068c4;
    assign coff[1934] = 256'h00001614ffff81ebffffe9ec00007e1500001614ffff81ebffffe9ec00007e15;
    assign coff[1935] = 256'hffff81ebffffe9ec00007e1500001614ffff81ebffffe9ec00007e1500001614;
    assign coff[1936] = 256'h00007f10fffff087ffff80f000000f7900007f10fffff087ffff80f000000f79;
    assign coff[1937] = 256'hfffff087ffff80f000000f7900007f10fffff087ffff80f000000f7900007f10;
    assign coff[1938] = 256'h00004ee8ffff9b36ffffb118000064ca00004ee8ffff9b36ffffb118000064ca;
    assign coff[1939] = 256'hffff9b36ffffb118000064ca00004ee8ffff9b36ffffb118000064ca00004ee8;
    assign coff[1940] = 256'h00006f78ffffc114ffff908800003eec00006f78ffffc114ffff908800003eec;
    assign coff[1941] = 256'hffffc114ffff908800003eec00006f78ffffc114ffff908800003eec00006f78;
    assign coff[1942] = 256'h00002254ffff84b0ffffddac00007b5000002254ffff84b0ffffddac00007b50;
    assign coff[1943] = 256'hffff84b0ffffddac00007b5000002254ffff84b0ffffddac00007b5000002254;
    assign coff[1944] = 256'h0000799affffd809ffff8666000027f70000799affffd809ffff8666000027f7;
    assign coff[1945] = 256'hffffd809ffff8666000027f70000799affffd809ffff8666000027f70000799a;
    assign coff[1946] = 256'h000039baffff8dc1ffffc6460000723f000039baffff8dc1ffffc6460000723f;
    assign coff[1947] = 256'hffff8dc1ffffc6460000723f000039baffff8dc1ffffc6460000723f000039ba;
    assign coff[1948] = 256'h0000610dffffac8bffff9ef3000053750000610dffffac8bffff9ef300005375;
    assign coff[1949] = 256'hffffac8bffff9ef3000053750000610dffffac8bffff9ef3000053750000610d;
    assign coff[1950] = 256'h0000099dffff805dfffff66300007fa30000099dffff805dfffff66300007fa3;
    assign coff[1951] = 256'hffff805dfffff66300007fa30000099dffff805dfffff66300007fa30000099d;
    assign coff[1952] = 256'h00007fabfffff6c8ffff80550000093800007fabfffff6c8ffff805500000938;
    assign coff[1953] = 256'hfffff6c8ffff80550000093800007fabfffff6c8ffff80550000093800007fab;
    assign coff[1954] = 256'h000053c1ffff9f35ffffac3f000060cb000053c1ffff9f35ffffac3f000060cb;
    assign coff[1955] = 256'hffff9f35ffffac3f000060cb000053c1ffff9f35ffffac3f000060cb000053c1;
    assign coff[1956] = 256'h0000726cffffc6a0ffff8d94000039600000726cffffc6a0ffff8d9400003960;
    assign coff[1957] = 256'hffffc6a0ffff8d94000039600000726cffffc6a0ffff8d94000039600000726c;
    assign coff[1958] = 256'h00002856ffff8686ffffd7aa0000797a00002856ffff8686ffffd7aa0000797a;
    assign coff[1959] = 256'hffff8686ffffd7aa0000797a00002856ffff8686ffffd7aa0000797a00002856;
    assign coff[1960] = 256'h00007b6affffde0dffff8496000021f300007b6affffde0dffff8496000021f3;
    assign coff[1961] = 256'hffffde0dffff8496000021f300007b6affffde0dffff8496000021f300007b6a;
    assign coff[1962] = 256'h00003f43ffff90baffffc0bd00006f4600003f43ffff90baffffc0bd00006f46;
    assign coff[1963] = 256'hffff90baffffc0bd00006f4600003f43ffff90baffffc0bd00006f4600003f43;
    assign coff[1964] = 256'h00006507ffffb168ffff9af900004e9800006507ffffb168ffff9af900004e98;
    assign coff[1965] = 256'hffffb168ffff9af900004e9800006507ffffb168ffff9af900004e9800006507;
    assign coff[1966] = 256'h00000fddffff80fdfffff02300007f0300000fddffff80fdfffff02300007f03;
    assign coff[1967] = 256'hffff80fdfffff02300007f0300000fddffff80fdfffff02300007f0300000fdd;
    assign coff[1968] = 256'h00007e26ffffea4fffff81da000015b100007e26ffffea4fffff81da000015b1;
    assign coff[1969] = 256'hffffea4fffff81da000015b100007e26ffffea4fffff81da000015b100007e26;
    assign coff[1970] = 256'h000049ddffff9776ffffb6230000688a000049ddffff9776ffffb6230000688a;
    assign coff[1971] = 256'hffff9776ffffb6230000688a000049ddffff9776ffffb6230000688a000049dd;
    assign coff[1972] = 256'h00006c3fffffbbb0ffff93c10000445000006c3fffffbbb0ffff93c100004450;
    assign coff[1973] = 256'hffffbbb0ffff93c10000445000006c3fffffbbb0ffff93c10000445000006c3f;
    assign coff[1974] = 256'h00001c3dffff8327ffffe3c300007cd900001c3dffff8327ffffe3c300007cd9;
    assign coff[1975] = 256'hffff8327ffffe3c300007cd900001c3dffff8327ffffe3c300007cd900001c3d;
    assign coff[1976] = 256'h0000777effffd21effff888200002de20000777effffd21effff888200002de2;
    assign coff[1977] = 256'hffffd21effff888200002de20000777effffd21effff888200002de20000777e;
    assign coff[1978] = 256'h0000340dffff8b10ffffcbf3000074f00000340dffff8b10ffffcbf3000074f0;
    assign coff[1979] = 256'hffff8b10ffffcbf3000074f00000340dffff8b10ffffcbf3000074f00000340d;
    assign coff[1980] = 256'h00005cd7ffffa7e2ffffa3290000581e00005cd7ffffa7e2ffffa3290000581e;
    assign coff[1981] = 256'hffffa7e2ffffa3290000581e00005cd7ffffa7e2ffffa3290000581e00005cd7;
    assign coff[1982] = 256'h00000356ffff800bfffffcaa00007ff500000356ffff800bfffffcaa00007ff5;
    assign coff[1983] = 256'hffff800bfffffcaa00007ff500000356ffff800bfffffcaa00007ff500000356;
    assign coff[1984] = 256'h00007fdbfffff9eaffff80250000061600007fdbfffff9eaffff802500000616;
    assign coff[1985] = 256'hfffff9eaffff80250000061600007fdbfffff9eaffff80250000061600007fdb;
    assign coff[1986] = 256'h0000561bffffa14affffa9e500005eb60000561bffffa14affffa9e500005eb6;
    assign coff[1987] = 256'hffffa14affffa9e500005eb60000561bffffa14affffa9e500005eb60000561b;
    assign coff[1988] = 256'h000073cbffffc973ffff8c350000368d000073cbffffc973ffff8c350000368d;
    assign coff[1989] = 256'hffffc973ffff8c350000368d000073cbffffc973ffff8c350000368d000073cb;
    assign coff[1990] = 256'h00002b4fffff878cffffd4b10000787400002b4fffff878cffffd4b100007874;
    assign coff[1991] = 256'hffff878cffffd4b10000787400002b4fffff878cffffd4b10000787400002b4f;
    assign coff[1992] = 256'h00007c36ffffe117ffff83ca00001ee900007c36ffffe117ffff83ca00001ee9;
    assign coff[1993] = 256'hffffe117ffff83ca00001ee900007c36ffffe117ffff83ca00001ee900007c36;
    assign coff[1994] = 256'h000041f9ffff9250ffffbe0700006db0000041f9ffff9250ffffbe0700006db0;
    assign coff[1995] = 256'hffff9250ffffbe0700006db0000041f9ffff9250ffffbe0700006db0000041f9;
    assign coff[1996] = 256'h000066edffffb3e9ffff991300004c17000066edffffb3e9ffff991300004c17;
    assign coff[1997] = 256'hffffb3e9ffff991300004c17000066edffffb3e9ffff991300004c17000066ed;
    assign coff[1998] = 256'h000012faffff816affffed0600007e96000012faffff816affffed0600007e96;
    assign coff[1999] = 256'hffff816affffed0600007e96000012faffff816affffed0600007e96000012fa;
    assign coff[2000] = 256'h00007ea5ffffed6affff815b0000129600007ea5ffffed6affff815b00001296;
    assign coff[2001] = 256'hffffed6affff815b0000129600007ea5ffffed6affff815b0000129600007ea5;
    assign coff[2002] = 256'h00004c68ffff994effffb398000066b200004c68ffff994effffb398000066b2;
    assign coff[2003] = 256'hffff994effffb398000066b200004c68ffff994effffb398000066b200004c68;
    assign coff[2004] = 256'h00006de4ffffbe5dffff921c000041a300006de4ffffbe5dffff921c000041a3;
    assign coff[2005] = 256'hffffbe5dffff921c000041a300006de4ffffbe5dffff921c000041a300006de4;
    assign coff[2006] = 256'h00001f4bffff83e2ffffe0b500007c1e00001f4bffff83e2ffffe0b500007c1e;
    assign coff[2007] = 256'hffff83e2ffffe0b500007c1e00001f4bffff83e2ffffe0b500007c1e00001f4b;
    assign coff[2008] = 256'h00007895ffffd510ffff876b00002af000007895ffffd510ffff876b00002af0;
    assign coff[2009] = 256'hffffd510ffff876b00002af000007895ffffd510ffff876b00002af000007895;
    assign coff[2010] = 256'h000036e8ffff8c60ffffc918000073a0000036e8ffff8c60ffffc918000073a0;
    assign coff[2011] = 256'hffff8c60ffffc918000073a0000036e8ffff8c60ffffc918000073a0000036e8;
    assign coff[2012] = 256'h00005ef9ffffaa30ffffa107000055d000005ef9ffffaa30ffffa107000055d0;
    assign coff[2013] = 256'hffffaa30ffffa107000055d000005ef9ffffaa30ffffa107000055d000005ef9;
    assign coff[2014] = 256'h0000067affff802afffff98600007fd60000067affff802afffff98600007fd6;
    assign coff[2015] = 256'hffff802afffff98600007fd60000067affff802afffff98600007fd60000067a;
    assign coff[2016] = 256'h00007f67fffff3a6ffff809900000c5a00007f67fffff3a6ffff809900000c5a;
    assign coff[2017] = 256'hfffff3a6ffff809900000c5a00007f67fffff3a6ffff809900000c5a00007f67;
    assign coff[2018] = 256'h0000515bffff9d2effffaea5000062d20000515bffff9d2effffaea5000062d2;
    assign coff[2019] = 256'hffff9d2effffaea5000062d20000515bffff9d2effffaea5000062d20000515b;
    assign coff[2020] = 256'h000070faffffc3d6ffff8f0600003c2a000070faffffc3d6ffff8f0600003c2a;
    assign coff[2021] = 256'hffffc3d6ffff8f0600003c2a000070faffffc3d6ffff8f0600003c2a000070fa;
    assign coff[2022] = 256'h00002558ffff8592ffffdaa800007a6e00002558ffff8592ffffdaa800007a6e;
    assign coff[2023] = 256'hffff8592ffffdaa800007a6e00002558ffff8592ffffdaa800007a6e00002558;
    assign coff[2024] = 256'h00007a8cffffdb08ffff8574000024f800007a8cffffdb08ffff8574000024f8;
    assign coff[2025] = 256'hffffdb08ffff8574000024f800007a8cffffdb08ffff8574000024f800007a8c;
    assign coff[2026] = 256'h00003c83ffff8f35ffffc37d000070cb00003c83ffff8f35ffffc37d000070cb;
    assign coff[2027] = 256'hffff8f35ffffc37d000070cb00003c83ffff8f35ffffc37d000070cb00003c83;
    assign coff[2028] = 256'h00006312ffffaef3ffff9cee0000510d00006312ffffaef3ffff9cee0000510d;
    assign coff[2029] = 256'hffffaef3ffff9cee0000510d00006312ffffaef3ffff9cee0000510d00006312;
    assign coff[2030] = 256'h00000cbeffff80a3fffff34200007f5d00000cbeffff80a3fffff34200007f5d;
    assign coff[2031] = 256'hffff80a3fffff34200007f5d00000cbeffff80a3fffff34200007f5d00000cbe;
    assign coff[2032] = 256'h00007d94ffffe739ffff826c000018c700007d94ffffe739ffff826c000018c7;
    assign coff[2033] = 256'hffffe739ffff826c000018c700007d94ffffe739ffff826c000018c700007d94;
    assign coff[2034] = 256'h00004747ffff95aeffffb8b900006a5200004747ffff95aeffffb8b900006a52;
    assign coff[2035] = 256'hffff95aeffffb8b900006a5200004747ffff95aeffffb8b900006a5200004747;
    assign coff[2036] = 256'h00006a89ffffb90dffff9577000046f300006a89ffffb90dffff9577000046f3;
    assign coff[2037] = 256'hffffb90dffff9577000046f300006a89ffffb90dffff9577000046f300006a89;
    assign coff[2038] = 256'h0000192affff827fffffe6d600007d810000192affff827fffffe6d600007d81;
    assign coff[2039] = 256'hffff827fffffe6d600007d810000192affff827fffffe6d600007d810000192a;
    assign coff[2040] = 256'h00007655ffffcf33ffff89ab000030cd00007655ffffcf33ffff89ab000030cd;
    assign coff[2041] = 256'hffffcf33ffff89ab000030cd00007655ffffcf33ffff89ab000030cd00007655;
    assign coff[2042] = 256'h0000312affff89d2ffffced60000762e0000312affff89d2ffffced60000762e;
    assign coff[2043] = 256'hffff89d2ffffced60000762e0000312affff89d2ffffced60000762e0000312a;
    assign coff[2044] = 256'h00005aa6ffffa5a1ffffa55a00005a5f00005aa6ffffa5a1ffffa55a00005a5f;
    assign coff[2045] = 256'hffffa5a1ffffa55a00005a5f00005aa6ffffa5a1ffffa55a00005a5f00005aa6;
    assign coff[2046] = 256'h00000032ffff8001ffffffce00007fff00000032ffff8001ffffffce00007fff;
    assign coff[2047] = 256'hffff8001ffffffce00007fff00000032ffff8001ffffffce00007fff00000032;

    always_ff @(posedge clk, negedge rst_n) begin
        if(~rst_n) begin
            data_o <= 'b0;
        end else if (valid == 1) begin
            data_o <= coff[addr_i];
        end else begin
            data_o <= 'b0;
        end
    end


endmodule