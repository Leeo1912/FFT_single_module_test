`timescale 1ns/1ps
module rom_recover_2n_twiddle
(
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic [13:0]              addr_i,
    output logic [63:0]              data_o
);

    logic [63:0] coff[8191:0];

    assign coff[0   ] = 64'h7fffffff00000000;
    assign coff[1   ] = 64'h5a82799aa57d8666;
    assign coff[2   ] = 64'h0000000080000000;
    assign coff[3   ] = 64'ha57d8666a57d8666;
    assign coff[4   ] = 64'h7641af3dcf043ab3;
    assign coff[5   ] = 64'h30fbc54d89be50c3;
    assign coff[6   ] = 64'hcf043ab389be50c3;
    assign coff[7   ] = 64'h89be50c3cf043ab3;
    assign coff[8   ] = 64'h7d8a5f40e70747c4;
    assign coff[9   ] = 64'h471cece79592675c;
    assign coff[10  ] = 64'he70747c48275a0c0;
    assign coff[11  ] = 64'h9592675cb8e31319;
    assign coff[12  ] = 64'h6a6d98a4b8e31319;
    assign coff[13  ] = 64'h18f8b83c8275a0c0;
    assign coff[14  ] = 64'hb8e313199592675c;
    assign coff[15  ] = 64'h8275a0c0e70747c4;
    assign coff[16  ] = 64'h70e2cbc6c3a94590;
    assign coff[17  ] = 64'h25280c5e8582faa5;
    assign coff[18  ] = 64'hc3a945908f1d343a;
    assign coff[19  ] = 64'h8582faa5dad7f3a2;
    assign coff[20  ] = 64'h7a7d055bdad7f3a2;
    assign coff[21  ] = 64'h3c56ba708f1d343a;
    assign coff[22  ] = 64'hdad7f3a28582faa5;
    assign coff[23  ] = 64'h8f1d343ac3a94590;
    assign coff[24  ] = 64'h7f62368ff3742ca2;
    assign coff[25  ] = 64'h5133cc949d0dfe54;
    assign coff[26  ] = 64'hf3742ca2809dc971;
    assign coff[27  ] = 64'h9d0dfe54aecc336c;
    assign coff[28  ] = 64'h62f201acaecc336c;
    assign coff[29  ] = 64'h0c8bd35e809dc971;
    assign coff[30  ] = 64'haecc336c9d0dfe54;
    assign coff[31  ] = 64'h809dc971f3742ca2;
    assign coff[32  ] = 64'h66cf8120b3c0200c;
    assign coff[33  ] = 64'h12c8106f8162aa04;
    assign coff[34  ] = 64'hb3c0200c99307ee0;
    assign coff[35  ] = 64'h8162aa04ed37ef91;
    assign coff[36  ] = 64'h7e9d55fced37ef91;
    assign coff[37  ] = 64'h4c3fdff499307ee0;
    assign coff[38  ] = 64'hed37ef918162aa04;
    assign coff[39  ] = 64'h99307ee0b3c0200c;
    assign coff[40  ] = 64'h7c29fbeee0e60685;
    assign coff[41  ] = 64'h41ce1e659235f2ec;
    assign coff[42  ] = 64'he0e6068583d60412;
    assign coff[43  ] = 64'h9235f2ecbe31e19b;
    assign coff[44  ] = 64'h6dca0d14be31e19b;
    assign coff[45  ] = 64'h1f19f97b83d60412;
    assign coff[46  ] = 64'hbe31e19b9235f2ec;
    assign coff[47  ] = 64'h83d60412e0e60685;
    assign coff[48  ] = 64'h73b5ebd1c945dfec;
    assign coff[49  ] = 64'h2b1f34eb877b7bec;
    assign coff[50  ] = 64'hc945dfec8c4a142f;
    assign coff[51  ] = 64'h877b7becd4e0cb15;
    assign coff[52  ] = 64'h78848414d4e0cb15;
    assign coff[53  ] = 64'h36ba20148c4a142f;
    assign coff[54  ] = 64'hd4e0cb15877b7bec;
    assign coff[55  ] = 64'h8c4a142fc945dfec;
    assign coff[56  ] = 64'h7fd8878ef9b82684;
    assign coff[57  ] = 64'h55f5a4d2a1288376;
    assign coff[58  ] = 64'hf9b8268480277872;
    assign coff[59  ] = 64'ha1288376aa0a5b2e;
    assign coff[60  ] = 64'h5ed77c8aaa0a5b2e;
    assign coff[61  ] = 64'h0647d97c80277872;
    assign coff[62  ] = 64'haa0a5b2ea1288376;
    assign coff[63  ] = 64'h80277872f9b82684;
    assign coff[64  ] = 64'h60ec3830ac64d510;
    assign coff[65  ] = 64'h096a90498058c94c;
    assign coff[66  ] = 64'hac64d5109f13c7d0;
    assign coff[67  ] = 64'h8058c94cf6956fb7;
    assign coff[68  ] = 64'h7fa736b4f6956fb7;
    assign coff[69  ] = 64'h539b2af09f13c7d0;
    assign coff[70  ] = 64'hf6956fb78058c94c;
    assign coff[71  ] = 64'h9f13c7d0ac64d510;
    assign coff[72  ] = 64'h798a23b1d7d946d8;
    assign coff[73  ] = 64'h398cdd328daad37b;
    assign coff[74  ] = 64'hd7d946d88675dc4f;
    assign coff[75  ] = 64'h8daad37bc67322ce;
    assign coff[76  ] = 64'h72552c85c67322ce;
    assign coff[77  ] = 64'h2826b9288675dc4f;
    assign coff[78  ] = 64'hc67322ce8daad37b;
    assign coff[79  ] = 64'h8675dc4fd7d946d8;
    assign coff[80  ] = 64'h6f5f02b2c0e8b648;
    assign coff[81  ] = 64'h2223a4c584a2fc62;
    assign coff[82  ] = 64'hc0e8b64890a0fd4e;
    assign coff[83  ] = 64'h84a2fc62dddc5b3b;
    assign coff[84  ] = 64'h7b5d039edddc5b3b;
    assign coff[85  ] = 64'h3f1749b890a0fd4e;
    assign coff[86  ] = 64'hdddc5b3b84a2fc62;
    assign coff[87  ] = 64'h90a0fd4ec0e8b648;
    assign coff[88  ] = 64'h7f0991c4f054d8d5;
    assign coff[89  ] = 64'h4ebfe8a59b1776da;
    assign coff[90  ] = 64'hf054d8d580f66e3c;
    assign coff[91  ] = 64'h9b1776dab140175b;
    assign coff[92  ] = 64'h64e88926b140175b;
    assign coff[93  ] = 64'h0fab272b80f66e3c;
    assign coff[94  ] = 64'hb140175b9b1776da;
    assign coff[95  ] = 64'h80f66e3cf054d8d5;
    assign coff[96  ] = 64'h68a69e81b64beacd;
    assign coff[97  ] = 64'h15e2144581e26c16;
    assign coff[98  ] = 64'hb64beacd9759617f;
    assign coff[99  ] = 64'h81e26c16ea1debbb;
    assign coff[100 ] = 64'h7e1d93eaea1debbb;
    assign coff[101 ] = 64'h49b415339759617f;
    assign coff[102 ] = 64'hea1debbb81e26c16;
    assign coff[103 ] = 64'h9759617fb64beacd;
    assign coff[104 ] = 64'h7ce3ceb2e3f47d96;
    assign coff[105 ] = 64'h447acd5093dbd6a0;
    assign coff[106 ] = 64'he3f47d96831c314e;
    assign coff[107 ] = 64'h93dbd6a0bb8532b0;
    assign coff[108 ] = 64'h6c242960bb8532b0;
    assign coff[109 ] = 64'h1c0b826a831c314e;
    assign coff[110 ] = 64'hbb8532b093dbd6a0;
    assign coff[111 ] = 64'h831c314ee3f47d96;
    assign coff[112 ] = 64'h7504d345cc210d79;
    assign coff[113 ] = 64'h2e110a628893b125;
    assign coff[114 ] = 64'hcc210d798afb2cbb;
    assign coff[115 ] = 64'h8893b125d1eef59e;
    assign coff[116 ] = 64'h776c4edbd1eef59e;
    assign coff[117 ] = 64'h33def2878afb2cbb;
    assign coff[118 ] = 64'hd1eef59e8893b125;
    assign coff[119 ] = 64'h8afb2cbbcc210d79;
    assign coff[120 ] = 64'h7ff62182fcdbd541;
    assign coff[121 ] = 64'h5842dd54a34bdf20;
    assign coff[122 ] = 64'hfcdbd5418009de7e;
    assign coff[123 ] = 64'ha34bdf20a7bd22ac;
    assign coff[124 ] = 64'h5cb420e0a7bd22ac;
    assign coff[125 ] = 64'h03242abf8009de7e;
    assign coff[126 ] = 64'ha7bd22aca34bdf20;
    assign coff[127 ] = 64'h8009de7efcdbd541;
    assign coff[128 ] = 64'h5dc79d7ca8e21106;
    assign coff[129 ] = 64'h04b6195d80163440;
    assign coff[130 ] = 64'ha8e21106a2386284;
    assign coff[131 ] = 64'h80163440fb49e6a3;
    assign coff[132 ] = 64'h7fe9cbc0fb49e6a3;
    assign coff[133 ] = 64'h571deefaa2386284;
    assign coff[134 ] = 64'hfb49e6a380163440;
    assign coff[135 ] = 64'ha2386284a8e21106;
    assign coff[136 ] = 64'h77fab989d3670446;
    assign coff[137 ] = 64'h354d90578ba0622f;
    assign coff[138 ] = 64'hd367044688054677;
    assign coff[139 ] = 64'h8ba0622fcab26fa9;
    assign coff[140 ] = 64'h745f9dd1cab26fa9;
    assign coff[141 ] = 64'h2c98fbba88054677;
    assign coff[142 ] = 64'hcab26fa98ba0622f;
    assign coff[143 ] = 64'h88054677d3670446;
    assign coff[144 ] = 64'h6cf934fcbcda3ecb;
    assign coff[145 ] = 64'h1d934fe58376b422;
    assign coff[146 ] = 64'hbcda3ecb9306cb04;
    assign coff[147 ] = 64'h8376b422e26cb01b;
    assign coff[148 ] = 64'h7c894bdee26cb01b;
    assign coff[149 ] = 64'h4325c1359306cb04;
    assign coff[150 ] = 64'he26cb01b8376b422;
    assign coff[151 ] = 64'h9306cb04bcda3ecb;
    assign coff[152 ] = 64'h7e5fe493ebaa894f;
    assign coff[153 ] = 64'h4afb6c989842f043;
    assign coff[154 ] = 64'hebaa894f81a01b6d;
    assign coff[155 ] = 64'h9842f043b5049368;
    assign coff[156 ] = 64'h67bd0fbdb5049368;
    assign coff[157 ] = 64'h145576b181a01b6d;
    assign coff[158 ] = 64'hb50493689842f043;
    assign coff[159 ] = 64'h81a01b6debaa894f;
    assign coff[160 ] = 64'h65ddfbd3b27e9d3c;
    assign coff[161 ] = 64'h1139f0cf812a1a3a;
    assign coff[162 ] = 64'hb27e9d3c9a22042d;
    assign coff[163 ] = 64'h812a1a3aeec60f31;
    assign coff[164 ] = 64'h7ed5e5c6eec60f31;
    assign coff[165 ] = 64'h4d8162c49a22042d;
    assign coff[166 ] = 64'heec60f31812a1a3a;
    assign coff[167 ] = 64'h9a22042db27e9d3c;
    assign coff[168 ] = 64'h7bc5e290df608fe4;
    assign coff[169 ] = 64'h4073f21d91695663;
    assign coff[170 ] = 64'hdf608fe4843a1d70;
    assign coff[171 ] = 64'h91695663bf8c0de3;
    assign coff[172 ] = 64'h6e96a99dbf8c0de3;
    assign coff[173 ] = 64'h209f701c843a1d70;
    assign coff[174 ] = 64'hbf8c0de391695663;
    assign coff[175 ] = 64'h843a1d70df608fe4;
    assign coff[176 ] = 64'h7307c3d0c7db6c50;
    assign coff[177 ] = 64'h29a3c48586f656d3;
    assign coff[178 ] = 64'hc7db6c508cf83c30;
    assign coff[179 ] = 64'h86f656d3d65c3b7b;
    assign coff[180 ] = 64'h7909a92dd65c3b7b;
    assign coff[181 ] = 64'h382493b08cf83c30;
    assign coff[182 ] = 64'hd65c3b7b86f656d3;
    assign coff[183 ] = 64'h8cf83c30c7db6c50;
    assign coff[184 ] = 64'h7fc25596f826a462;
    assign coff[185 ] = 64'h54ca0a4ba01c4c73;
    assign coff[186 ] = 64'hf826a462803daa6a;
    assign coff[187 ] = 64'ha01c4c73ab35f5b5;
    assign coff[188 ] = 64'h5fe3b38dab35f5b5;
    assign coff[189 ] = 64'h07d95b9e803daa6a;
    assign coff[190 ] = 64'hab35f5b5a01c4c73;
    assign coff[191 ] = 64'h803daa6af826a462;
    assign coff[192 ] = 64'h61f1003fad96ed92;
    assign coff[193 ] = 64'h0afb68058078d40d;
    assign coff[194 ] = 64'had96ed929e0effc1;
    assign coff[195 ] = 64'h8078d40df50497fb;
    assign coff[196 ] = 64'h7f872bf3f50497fb;
    assign coff[197 ] = 64'h5269126e9e0effc1;
    assign coff[198 ] = 64'hf50497fb8078d40d;
    assign coff[199 ] = 64'h9e0effc1ad96ed92;
    assign coff[200 ] = 64'h7a05eeadd957de7a;
    assign coff[201 ] = 64'h3af2eeb78e61d32e;
    assign coff[202 ] = 64'hd957de7a85fa1153;
    assign coff[203 ] = 64'h8e61d32ec50d1149;
    assign coff[204 ] = 64'h719e2cd2c50d1149;
    assign coff[205 ] = 64'h26a8218685fa1153;
    assign coff[206 ] = 64'hc50d11498e61d32e;
    assign coff[207 ] = 64'h85fa1153d957de7a;
    assign coff[208 ] = 64'h7023109ac247cd5a;
    assign coff[209 ] = 64'h23a6887f85109cdd;
    assign coff[210 ] = 64'hc247cd5a8fdcef66;
    assign coff[211 ] = 64'h85109cdddc597781;
    assign coff[212 ] = 64'h7aef6323dc597781;
    assign coff[213 ] = 64'h3db832a68fdcef66;
    assign coff[214 ] = 64'hdc59778185109cdd;
    assign coff[215 ] = 64'h8fdcef66c247cd5a;
    assign coff[216 ] = 64'h7f3857f6f1e43d1c;
    assign coff[217 ] = 64'h4ffb654d9c10cd70;
    assign coff[218 ] = 64'hf1e43d1c80c7a80a;
    assign coff[219 ] = 64'h9c10cd70b0049ab3;
    assign coff[220 ] = 64'h63ef3290b0049ab3;
    assign coff[221 ] = 64'h0e1bc2e480c7a80a;
    assign coff[222 ] = 64'hb0049ab39c10cd70;
    assign coff[223 ] = 64'h80c7a80af1e43d1c;
    assign coff[224 ] = 64'h698c246cb796199b;
    assign coff[225 ] = 64'h176dd9de82299971;
    assign coff[226 ] = 64'hb796199b9673db94;
    assign coff[227 ] = 64'h82299971e8922622;
    assign coff[228 ] = 64'h7dd6668fe8922622;
    assign coff[229 ] = 64'h4869e6659673db94;
    assign coff[230 ] = 64'he892262282299971;
    assign coff[231 ] = 64'h9673db94b796199b;
    assign coff[232 ] = 64'h7d3980ece57d5fda;
    assign coff[233 ] = 64'h45cd358f94b50d87;
    assign coff[234 ] = 64'he57d5fda82c67f14;
    assign coff[235 ] = 64'h94b50d87ba32ca71;
    assign coff[236 ] = 64'h6b4af279ba32ca71;
    assign coff[237 ] = 64'h1a82a02682c67f14;
    assign coff[238 ] = 64'hba32ca7194b50d87;
    assign coff[239 ] = 64'h82c67f14e57d5fda;
    assign coff[240 ] = 64'h75a585cfcd91ab39;
    assign coff[241 ] = 64'h2f8752628926b677;
    assign coff[242 ] = 64'hcd91ab398a5a7a31;
    assign coff[243 ] = 64'h8926b677d078ad9e;
    assign coff[244 ] = 64'h76d94989d078ad9e;
    assign coff[245 ] = 64'h326e54c78a5a7a31;
    assign coff[246 ] = 64'hd078ad9e8926b677;
    assign coff[247 ] = 64'h8a5a7a31cd91ab39;
    assign coff[248 ] = 64'h7ffd885afe6de2e0;
    assign coff[249 ] = 64'h59646498a462eeac;
    assign coff[250 ] = 64'hfe6de2e0800277a6;
    assign coff[251 ] = 64'ha462eeaca69b9b68;
    assign coff[252 ] = 64'h5b9d1154a69b9b68;
    assign coff[253 ] = 64'h01921d20800277a6;
    assign coff[254 ] = 64'ha69b9b68a462eeac;
    assign coff[255 ] = 64'h800277a6fe6de2e0;
    assign coff[256 ] = 64'h5c290acca72bf174;
    assign coff[257 ] = 64'h025b26d780058d2f;
    assign coff[258 ] = 64'ha72bf174a3d6f534;
    assign coff[259 ] = 64'h80058d2ffda4d929;
    assign coff[260 ] = 64'h7ffa72d1fda4d929;
    assign coff[261 ] = 64'h58d40e8ca3d6f534;
    assign coff[262 ] = 64'hfda4d92980058d2f;
    assign coff[263 ] = 64'ha3d6f534a72bf174;
    assign coff[264 ] = 64'h77235f2dd13397e2;
    assign coff[265 ] = 64'h3326e2c38aaa42b4;
    assign coff[266 ] = 64'hd13397e288dca0d3;
    assign coff[267 ] = 64'h8aaa42b4ccd91d3d;
    assign coff[268 ] = 64'h7555bd4cccd91d3d;
    assign coff[269 ] = 64'h2ecc681e88dca0d3;
    assign coff[270 ] = 64'hccd91d3d8aaa42b4;
    assign coff[271 ] = 64'h88dca0d3d13397e2;
    assign coff[272 ] = 64'h6bb812d1badba943;
    assign coff[273 ] = 64'h1b4732ef82f0bde8;
    assign coff[274 ] = 64'hbadba9439447ed2f;
    assign coff[275 ] = 64'h82f0bde8e4b8cd11;
    assign coff[276 ] = 64'h7d0f4218e4b8cd11;
    assign coff[277 ] = 64'h452456bd9447ed2f;
    assign coff[278 ] = 64'he4b8cd1182f0bde8;
    assign coff[279 ] = 64'h9447ed2fbadba943;
    assign coff[280 ] = 64'h7dfa98a8e957ecfb;
    assign coff[281 ] = 64'h490f57ee96e61ce0;
    assign coff[282 ] = 64'he957ecfb82056758;
    assign coff[283 ] = 64'h96e61ce0b6f0a812;
    assign coff[284 ] = 64'h6919e320b6f0a812;
    assign coff[285 ] = 64'h16a8130582056758;
    assign coff[286 ] = 64'hb6f0a81296e61ce0;
    assign coff[287 ] = 64'h82056758e957ecfb;
    assign coff[288 ] = 64'h646c59bfb0a1f71d;
    assign coff[289 ] = 64'h0ee3876680de6e4c;
    assign coff[290 ] = 64'hb0a1f71d9b93a641;
    assign coff[291 ] = 64'h80de6e4cf11c789a;
    assign coff[292 ] = 64'h7f2191b4f11c789a;
    assign coff[293 ] = 64'h4f5e08e39b93a641;
    assign coff[294 ] = 64'hf11c789a80de6e4c;
    assign coff[295 ] = 64'h9b93a641b0a1f71d;
    assign coff[296 ] = 64'h7b26cb4fdd1abe51;
    assign coff[297 ] = 64'h3e680b2c903e6c7b;
    assign coff[298 ] = 64'hdd1abe5184d934b1;
    assign coff[299 ] = 64'h903e6c7bc197f4d4;
    assign coff[300 ] = 64'h6fc19385c197f4d4;
    assign coff[301 ] = 64'h22e541af84d934b1;
    assign coff[302 ] = 64'hc197f4d4903e6c7b;
    assign coff[303 ] = 64'h84d934b1dd1abe51;
    assign coff[304 ] = 64'h71fa3949c5bfd22e;
    assign coff[305 ] = 64'h27679df486376092;
    assign coff[306 ] = 64'hc5bfd22e8e05c6b7;
    assign coff[307 ] = 64'h86376092d898620c;
    assign coff[308 ] = 64'h79c89f6ed898620c;
    assign coff[309 ] = 64'h3a402dd28e05c6b7;
    assign coff[310 ] = 64'hd898620c86376092;
    assign coff[311 ] = 64'h8e05c6b7c5bfd22e;
    assign coff[312 ] = 64'h7f97cebdf5ccf743;
    assign coff[313 ] = 64'h530285189e90eb94;
    assign coff[314 ] = 64'hf5ccf74380683143;
    assign coff[315 ] = 64'h9e90eb94acfd7ae8;
    assign coff[316 ] = 64'h616f146cacfd7ae8;
    assign coff[317 ] = 64'h0a3308bd80683143;
    assign coff[318 ] = 64'hacfd7ae89e90eb94;
    assign coff[319 ] = 64'h80683143f5ccf743;
    assign coff[320 ] = 64'h60686ccfabccfd83;
    assign coff[321 ] = 64'h08a2009a804a9c4d;
    assign coff[322 ] = 64'habccfd839f979331;
    assign coff[323 ] = 64'h804a9c4df75dff66;
    assign coff[324 ] = 64'h7fb563b3f75dff66;
    assign coff[325 ] = 64'h5433027d9f979331;
    assign coff[326 ] = 64'hf75dff66804a9c4d;
    assign coff[327 ] = 64'h9f979331abccfd83;
    assign coff[328 ] = 64'h794a7c12d71a8eb5;
    assign coff[329 ] = 64'h38d8fe938d50fa59;
    assign coff[330 ] = 64'hd71a8eb586b583ee;
    assign coff[331 ] = 64'h8d50fa59c727016d;
    assign coff[332 ] = 64'h72af05a7c727016d;
    assign coff[333 ] = 64'h28e5714b86b583ee;
    assign coff[334 ] = 64'hc727016d8d50fa59;
    assign coff[335 ] = 64'h86b583eed71a8eb5;
    assign coff[336 ] = 64'h6efb5f12c03a1368;
    assign coff[337 ] = 64'h2161b3a0846df477;
    assign coff[338 ] = 64'hc03a13689104a0ee;
    assign coff[339 ] = 64'h846df477de9e4c60;
    assign coff[340 ] = 64'h7b920b89de9e4c60;
    assign coff[341 ] = 64'h3fc5ec989104a0ee;
    assign coff[342 ] = 64'hde9e4c60846df477;
    assign coff[343 ] = 64'h9104a0eec03a1368;
    assign coff[344 ] = 64'h7ef05860ef8d5fb8;
    assign coff[345 ] = 64'h4e2106179a9c406e;
    assign coff[346 ] = 64'hef8d5fb8810fa7a0;
    assign coff[347 ] = 64'h9a9c406eb1def9e9;
    assign coff[348 ] = 64'h6563bf92b1def9e9;
    assign coff[349 ] = 64'h1072a048810fa7a0;
    assign coff[350 ] = 64'hb1def9e99a9c406e;
    assign coff[351 ] = 64'h810fa7a0ef8d5fb8;
    assign coff[352 ] = 64'h683257abb5a7e362;
    assign coff[353 ] = 64'h151bdf8681c0a801;
    assign coff[354 ] = 64'hb5a7e36297cda855;
    assign coff[355 ] = 64'h81c0a801eae4207a;
    assign coff[356 ] = 64'h7e3f57ffeae4207a;
    assign coff[357 ] = 64'h4a581c9e97cda855;
    assign coff[358 ] = 64'heae4207a81c0a801;
    assign coff[359 ] = 64'h97cda855b5a7e362;
    assign coff[360 ] = 64'h7cb72724e330734d;
    assign coff[361 ] = 64'h43d09aed9370cae4;
    assign coff[362 ] = 64'he330734d8348d8dc;
    assign coff[363 ] = 64'h9370cae4bc2f6513;
    assign coff[364 ] = 64'h6c8f351cbc2f6513;
    assign coff[365 ] = 64'h1ccf8cb38348d8dc;
    assign coff[366 ] = 64'hbc2f65139370cae4;
    assign coff[367 ] = 64'h8348d8dce330734d;
    assign coff[368 ] = 64'h74b2c884cb697db0;
    assign coff[369 ] = 64'h2d553afc884be821;
    assign coff[370 ] = 64'hcb697db08b4d377c;
    assign coff[371 ] = 64'h884be821d2aac504;
    assign coff[372 ] = 64'h77b417dfd2aac504;
    assign coff[373 ] = 64'h349682508b4d377c;
    assign coff[374 ] = 64'hd2aac504884be821;
    assign coff[375 ] = 64'h8b4d377ccb697db0;
    assign coff[376 ] = 64'h7ff09478fc12d91a;
    assign coff[377 ] = 64'h57b0d256a2c1adc9;
    assign coff[378 ] = 64'hfc12d91a800f6b88;
    assign coff[379 ] = 64'ha2c1adc9a84f2daa;
    assign coff[380 ] = 64'h5d3e5237a84f2daa;
    assign coff[381 ] = 64'h03ed26e6800f6b88;
    assign coff[382 ] = 64'ha84f2daaa2c1adc9;
    assign coff[383 ] = 64'h800f6b88fc12d91a;
    assign coff[384 ] = 64'h5e50015da975cb57;
    assign coff[385 ] = 64'h057f0035801e3895;
    assign coff[386 ] = 64'ha975cb57a1affea3;
    assign coff[387 ] = 64'h801e3895fa80ffcb;
    assign coff[388 ] = 64'h7fe1c76bfa80ffcb;
    assign coff[389 ] = 64'h568a34a9a1affea3;
    assign coff[390 ] = 64'hfa80ffcb801e3895;
    assign coff[391 ] = 64'ha1affea3a975cb57;
    assign coff[392 ] = 64'h78403329d423b191;
    assign coff[393 ] = 64'h36041ad98bf4ac05;
    assign coff[394 ] = 64'hd423b19187bfccd7;
    assign coff[395 ] = 64'h8bf4ac05c9fbe527;
    assign coff[396 ] = 64'h740b53fbc9fbe527;
    assign coff[397 ] = 64'h2bdc4e6f87bfccd7;
    assign coff[398 ] = 64'hc9fbe5278bf4ac05;
    assign coff[399 ] = 64'h87bfccd7d423b191;
    assign coff[400 ] = 64'h6d6227fabd85be30;
    assign coff[401 ] = 64'h1e56ca1e83a5c2b0;
    assign coff[402 ] = 64'hbd85be30929dd806;
    assign coff[403 ] = 64'h83a5c2b0e1a935e2;
    assign coff[404 ] = 64'h7c5a3d50e1a935e2;
    assign coff[405 ] = 64'h427a41d0929dd806;
    assign coff[406 ] = 64'he1a935e283a5c2b0;
    assign coff[407 ] = 64'h929dd806bd85be30;
    assign coff[408 ] = 64'h7e7f3957ec71244f;
    assign coff[409 ] = 64'h4b9e039098b93828;
    assign coff[410 ] = 64'hec71244f8180c6a9;
    assign coff[411 ] = 64'h98b93828b461fc70;
    assign coff[412 ] = 64'h6746c7d8b461fc70;
    assign coff[413 ] = 64'h138edbb18180c6a9;
    assign coff[414 ] = 64'hb461fc7098b93828;
    assign coff[415 ] = 64'h8180c6a9ec71244f;
    assign coff[416 ] = 64'h66573cbbb31effcc;
    assign coff[417 ] = 64'h120116d58145c5c7;
    assign coff[418 ] = 64'hb31effcc99a8c345;
    assign coff[419 ] = 64'h8145c5c7edfee92b;
    assign coff[420 ] = 64'h7eba3a39edfee92b;
    assign coff[421 ] = 64'h4ce1003499a8c345;
    assign coff[422 ] = 64'hedfee92b8145c5c7;
    assign coff[423 ] = 64'h99a8c345b31effcc;
    assign coff[424 ] = 64'h7bf88830e02323e5;
    assign coff[425 ] = 64'h4121589b91cf1cb6;
    assign coff[426 ] = 64'he02323e5840777d0;
    assign coff[427 ] = 64'h91cf1cb6bedea765;
    assign coff[428 ] = 64'h6e30e34abedea765;
    assign coff[429 ] = 64'h1fdcdc1b840777d0;
    assign coff[430 ] = 64'hbedea76591cf1cb6;
    assign coff[431 ] = 64'h840777d0e02323e5;
    assign coff[432 ] = 64'h735f6626c89061ba;
    assign coff[433 ] = 64'h2a61b1018738545e;
    assign coff[434 ] = 64'hc89061ba8ca099da;
    assign coff[435 ] = 64'h8738545ed59e4eff;
    assign coff[436 ] = 64'h78c7aba2d59e4eff;
    assign coff[437 ] = 64'h376f9e468ca099da;
    assign coff[438 ] = 64'hd59e4eff8738545e;
    assign coff[439 ] = 64'h8ca099dac89061ba;
    assign coff[440 ] = 64'h7fce0c3ef8ef5cbb;
    assign coff[441 ] = 64'h556040e2a0a1f24d;
    assign coff[442 ] = 64'hf8ef5cbb8031f3c2;
    assign coff[443 ] = 64'ha0a1f24daa9fbf1e;
    assign coff[444 ] = 64'h5f5e0db3aa9fbf1e;
    assign coff[445 ] = 64'h0710a3458031f3c2;
    assign coff[446 ] = 64'haa9fbf1ea0a1f24d;
    assign coff[447 ] = 64'h8031f3c2f8ef5cbb;
    assign coff[448 ] = 64'h6271fa69ae312b92;
    assign coff[449 ] = 64'h0bc3ac35808ab180;
    assign coff[450 ] = 64'hae312b929d8e0597;
    assign coff[451 ] = 64'h808ab180f43c53cb;
    assign coff[452 ] = 64'h7f754e80f43c53cb;
    assign coff[453 ] = 64'h51ced46e9d8e0597;
    assign coff[454 ] = 64'hf43c53cb808ab180;
    assign coff[455 ] = 64'h9d8e0597ae312b92;
    assign coff[456 ] = 64'h7a4210d8da17ba4a;
    assign coff[457 ] = 64'h3ba51e298ebef7fb;
    assign coff[458 ] = 64'hda17ba4a85bdef28;
    assign coff[459 ] = 64'h8ebef7fbc45ae1d7;
    assign coff[460 ] = 64'h71410805c45ae1d7;
    assign coff[461 ] = 64'h25e845b685bdef28;
    assign coff[462 ] = 64'hc45ae1d78ebef7fb;
    assign coff[463 ] = 64'h85bdef28da17ba4a;
    assign coff[464 ] = 64'h708378ffc2f83e2a;
    assign coff[465 ] = 64'h246777588549345c;
    assign coff[466 ] = 64'hc2f83e2a8f7c8701;
    assign coff[467 ] = 64'h8549345cdb9888a8;
    assign coff[468 ] = 64'h7ab6cba4db9888a8;
    assign coff[469 ] = 64'h3d07c1d68f7c8701;
    assign coff[470 ] = 64'hdb9888a88549345c;
    assign coff[471 ] = 64'h8f7c8701c2f83e2a;
    assign coff[472 ] = 64'h7f4de451f2ac246e;
    assign coff[473 ] = 64'h5097fc5e9c8eeb34;
    assign coff[474 ] = 64'hf2ac246e80b21baf;
    assign coff[475 ] = 64'h9c8eeb34af6803a2;
    assign coff[476 ] = 64'h637114ccaf6803a2;
    assign coff[477 ] = 64'h0d53db9280b21baf;
    assign coff[478 ] = 64'haf6803a29c8eeb34;
    assign coff[479 ] = 64'h80b21baff2ac246e;
    assign coff[480 ] = 64'h69fd614ab83c3dd1;
    assign coff[481 ] = 64'h183366e9824f0208;
    assign coff[482 ] = 64'hb83c3dd196029eb6;
    assign coff[483 ] = 64'h824f0208e7cc9917;
    assign coff[484 ] = 64'h7db0fdf8e7cc9917;
    assign coff[485 ] = 64'h47c3c22f96029eb6;
    assign coff[486 ] = 64'he7cc9917824f0208;
    assign coff[487 ] = 64'h96029eb6b83c3dd1;
    assign coff[488 ] = 64'h7d628ac6e642340d;
    assign coff[489 ] = 64'h467568289523369c;
    assign coff[490 ] = 64'he642340d829d753a;
    assign coff[491 ] = 64'h9523369cb98a97d8;
    assign coff[492 ] = 64'h6adcc964b98a97d8;
    assign coff[493 ] = 64'h19bdcbf3829d753a;
    assign coff[494 ] = 64'hb98a97d89523369c;
    assign coff[495 ] = 64'h829d753ae642340d;
    assign coff[496 ] = 64'h75f42c0bce4ab5a2;
    assign coff[497 ] = 64'h3041c7618971f15a;
    assign coff[498 ] = 64'hce4ab5a28a0bd3f5;
    assign coff[499 ] = 64'h8971f15acfbe389f;
    assign coff[500 ] = 64'h768e0ea6cfbe389f;
    assign coff[501 ] = 64'h31b54a5e8a0bd3f5;
    assign coff[502 ] = 64'hcfbe389f8971f15a;
    assign coff[503 ] = 64'h8a0bd3f5ce4ab5a2;
    assign coff[504 ] = 64'h7fff6216ff36f078;
    assign coff[505 ] = 64'h59f3de12a4efca31;
    assign coff[506 ] = 64'hff36f07880009dea;
    assign coff[507 ] = 64'ha4efca31a60c21ee;
    assign coff[508 ] = 64'h5b1035cfa60c21ee;
    assign coff[509 ] = 64'h00c90f8880009dea;
    assign coff[510 ] = 64'ha60c21eea4efca31;
    assign coff[511 ] = 64'h80009deaff36f078;
    assign coff[512 ] = 64'h5b56bfbda653c303;
    assign coff[513 ] = 64'h012d96b18001634e;
    assign coff[514 ] = 64'ha653c303a4a94043;
    assign coff[515 ] = 64'h8001634efed2694f;
    assign coff[516 ] = 64'h7ffe9cb2fed2694f;
    assign coff[517 ] = 64'h59ac3cfda4a94043;
    assign coff[518 ] = 64'hfed2694f8001634e;
    assign coff[519 ] = 64'ha4a94043a653c303;
    assign coff[520 ] = 64'h76b3d0b4d01b6459;
    assign coff[521 ] = 64'h3211df048a3302be;
    assign coff[522 ] = 64'hd01b6459894c2f4c;
    assign coff[523 ] = 64'h8a3302becdee20fc;
    assign coff[524 ] = 64'h75ccfd42cdee20fc;
    assign coff[525 ] = 64'h2fe49ba7894c2f4c;
    assign coff[526 ] = 64'hcdee20fc8a3302be;
    assign coff[527 ] = 64'h894c2f4cd01b6459;
    assign coff[528 ] = 64'h6b13fef5b9de9b83;
    assign coff[529 ] = 64'h1a203e1b82b1d381;
    assign coff[530 ] = 64'hb9de9b8394ec010b;
    assign coff[531 ] = 64'h82b1d381e5dfc1e5;
    assign coff[532 ] = 64'h7d4e2c7fe5dfc1e5;
    assign coff[533 ] = 64'h4621647d94ec010b;
    assign coff[534 ] = 64'he5dfc1e582b1d381;
    assign coff[535 ] = 64'h94ec010bb9de9b83;
    assign coff[536 ] = 64'h7dc3d90de82f5844;
    assign coff[537 ] = 64'h4816ea86963b1c86;
    assign coff[538 ] = 64'he82f5844823c26f3;
    assign coff[539 ] = 64'h963b1c86b7e9157a;
    assign coff[540 ] = 64'h69c4e37ab7e9157a;
    assign coff[541 ] = 64'h17d0a7bc823c26f3;
    assign coff[542 ] = 64'hb7e9157a963b1c86;
    assign coff[543 ] = 64'h823c26f3e82f5844;
    assign coff[544 ] = 64'h63b0426dafb63667;
    assign coff[545 ] = 64'h0db7d37680bcba9d;
    assign coff[546 ] = 64'hafb636679c4fbd93;
    assign coff[547 ] = 64'h80bcba9df2482c8a;
    assign coff[548 ] = 64'h7f434563f2482c8a;
    assign coff[549 ] = 64'h5049c9999c4fbd93;
    assign coff[550 ] = 64'hf2482c8a80bcba9d;
    assign coff[551 ] = 64'h9c4fbd93afb63667;
    assign coff[552 ] = 64'h7ad33d45dbf8f4f8;
    assign coff[553 ] = 64'h3d600d2c8fac988f;
    assign coff[554 ] = 64'hdbf8f4f8852cc2bb;
    assign coff[555 ] = 64'h8fac988fc29ff2d4;
    assign coff[556 ] = 64'h70536771c29ff2d4;
    assign coff[557 ] = 64'h24070b08852cc2bb;
    assign coff[558 ] = 64'hc29ff2d48fac988f;
    assign coff[559 ] = 64'h852cc2bbdbf8f4f8;
    assign coff[560 ] = 64'h716fbd68c4b3e746;
    assign coff[561 ] = 64'h26483f6c85dbda91;
    assign coff[562 ] = 64'hc4b3e7468e904298;
    assign coff[563 ] = 64'h85dbda91d9b7c094;
    assign coff[564 ] = 64'h7a24256fd9b7c094;
    assign coff[565 ] = 64'h3b4c18ba8e904298;
    assign coff[566 ] = 64'hd9b7c09485dbda91;
    assign coff[567 ] = 64'h8e904298c4b3e746;
    assign coff[568 ] = 64'h7f7e648cf4a07261;
    assign coff[569 ] = 64'h521c0cc29dce6463;
    assign coff[570 ] = 64'hf4a0726180819b74;
    assign coff[571 ] = 64'h9dce6463ade3f33e;
    assign coff[572 ] = 64'h62319b9dade3f33e;
    assign coff[573 ] = 64'h0b5f8d9f80819b74;
    assign coff[574 ] = 64'hade3f33e9dce6463;
    assign coff[575 ] = 64'h80819b74f4a07261;
    assign coff[576 ] = 64'h5fa0fe1faaeac02c;
    assign coff[577 ] = 64'h077501be8037a7ac;
    assign coff[578 ] = 64'haaeac02ca05f01e1;
    assign coff[579 ] = 64'h8037a7acf88afe42;
    assign coff[580 ] = 64'h7fc85854f88afe42;
    assign coff[581 ] = 64'h55153fd4a05f01e1;
    assign coff[582 ] = 64'hf88afe428037a7ac;
    assign coff[583 ] = 64'ha05f01e1aaeac02c;
    assign coff[584 ] = 64'h78e8cfb2d5fd3848;
    assign coff[585 ] = 64'h37ca2a308ccc477d;
    assign coff[586 ] = 64'hd5fd38488717304e;
    assign coff[587 ] = 64'h8ccc477dc835d5d0;
    assign coff[588 ] = 64'h7333b883c835d5d0;
    assign coff[589 ] = 64'h2a02c7b88717304e;
    assign coff[590 ] = 64'hc835d5d08ccc477d;
    assign coff[591 ] = 64'h8717304ed5fd3848;
    assign coff[592 ] = 64'h6e63e87fbf3546a8;
    assign coff[593 ] = 64'h203e300d8420a46c;
    assign coff[594 ] = 64'hbf3546a8919c1781;
    assign coff[595 ] = 64'h8420a46cdfc1cff3;
    assign coff[596 ] = 64'h7bdf5b94dfc1cff3;
    assign coff[597 ] = 64'h40cab958919c1781;
    assign coff[598 ] = 64'hdfc1cff38420a46c;
    assign coff[599 ] = 64'h919c1781bf3546a8;
    assign coff[600 ] = 64'h7ec8371aee6276bf;
    assign coff[601 ] = 64'h4d31494b99e5443b;
    assign coff[602 ] = 64'hee6276bf8137c8e6;
    assign coff[603 ] = 64'h99e5443bb2ceb6b5;
    assign coff[604 ] = 64'h661abbc5b2ceb6b5;
    assign coff[605 ] = 64'h119d89418137c8e6;
    assign coff[606 ] = 64'hb2ceb6b599e5443b;
    assign coff[607 ] = 64'h8137c8e6ee6276bf;
    assign coff[608 ] = 64'h67820bb7b4b330b3;
    assign coff[609 ] = 64'h13f22f5881904a0c;
    assign coff[610 ] = 64'hb4b330b3987df449;
    assign coff[611 ] = 64'h81904a0cec0dd0a8;
    assign coff[612 ] = 64'h7e6fb5f4ec0dd0a8;
    assign coff[613 ] = 64'h4b4ccf4d987df449;
    assign coff[614 ] = 64'hec0dd0a881904a0c;
    assign coff[615 ] = 64'h987df449b4b330b3;
    assign coff[616 ] = 64'h7c71eaf9e20ae9c1;
    assign coff[617 ] = 64'h42d0161e92d22fd9;
    assign coff[618 ] = 64'he20ae9c1838e1507;
    assign coff[619 ] = 64'h92d22fd9bd2fe9e2;
    assign coff[620 ] = 64'h6d2dd027bd2fe9e2;
    assign coff[621 ] = 64'h1df5163f838e1507;
    assign coff[622 ] = 64'hbd2fe9e292d22fd9;
    assign coff[623 ] = 64'h838e1507e20ae9c1;
    assign coff[624 ] = 64'h74359cbdca5719db;
    assign coff[625 ] = 64'h2c3ab2b987e2649b;
    assign coff[626 ] = 64'hca5719db8bca6343;
    assign coff[627 ] = 64'h87e2649bd3c54d47;
    assign coff[628 ] = 64'h781d9b65d3c54d47;
    assign coff[629 ] = 64'h35a8e6258bca6343;
    assign coff[630 ] = 64'hd3c54d4787e2649b;
    assign coff[631 ] = 64'h8bca6343ca5719db;
    assign coff[632 ] = 64'h7fe5f108fae571a4;
    assign coff[633 ] = 64'h56d42c99a1f41392;
    assign coff[634 ] = 64'hfae571a4801a0ef8;
    assign coff[635 ] = 64'ha1f41392a92bd367;
    assign coff[636 ] = 64'h5e0bec6ea92bd367;
    assign coff[637 ] = 64'h051a8e5c801a0ef8;
    assign coff[638 ] = 64'ha92bd367a1f41392;
    assign coff[639 ] = 64'h801a0ef8fae571a4;
    assign coff[640 ] = 64'h5d8314b1a8988463;
    assign coff[641 ] = 64'h0451a1778012a86f;
    assign coff[642 ] = 64'ha8988463a27ceb4f;
    assign coff[643 ] = 64'h8012a86ffbae5e89;
    assign coff[644 ] = 64'h7fed5791fbae5e89;
    assign coff[645 ] = 64'h57677b9da27ceb4f;
    assign coff[646 ] = 64'hfbae5e898012a86f;
    assign coff[647 ] = 64'ha27ceb4fa8988463;
    assign coff[648 ] = 64'h77d78daad308d6c7;
    assign coff[649 ] = 64'h34f219a88b76a8e4;
    assign coff[650 ] = 64'hd308d6c788287256;
    assign coff[651 ] = 64'h8b76a8e4cb0de658;
    assign coff[652 ] = 64'h7489571ccb0de658;
    assign coff[653 ] = 64'h2cf7293988287256;
    assign coff[654 ] = 64'hcb0de6588b76a8e4;
    assign coff[655 ] = 64'h88287256d308d6c7;
    assign coff[656 ] = 64'h6cc45698bc84bd1f;
    assign coff[657 ] = 64'h1d31774d835fa00f;
    assign coff[658 ] = 64'hbc84bd1f933ba968;
    assign coff[659 ] = 64'h835fa00fe2ce88b3;
    assign coff[660 ] = 64'h7ca05ff1e2ce88b3;
    assign coff[661 ] = 64'h437b42e1933ba968;
    assign coff[662 ] = 64'he2ce88b3835fa00f;
    assign coff[663 ] = 64'h933ba968bc84bd1f;
    assign coff[664 ] = 64'h7e4fc53eeb474e81;
    assign coff[665 ] = 64'h4aa9dba298082c3b;
    assign coff[666 ] = 64'heb474e8181b03ac2;
    assign coff[667 ] = 64'h98082c3bb556245e;
    assign coff[668 ] = 64'h67f7d3c5b556245e;
    assign coff[669 ] = 64'h14b8b17f81b03ac2;
    assign coff[670 ] = 64'hb556245e98082c3b;
    assign coff[671 ] = 64'h81b03ac2eb474e81;
    assign coff[672 ] = 64'h65a0fd0bb22eb392;
    assign coff[673 ] = 64'h10d64dbd811cb9ca;
    assign coff[674 ] = 64'hb22eb3929a5f02f5;
    assign coff[675 ] = 64'h811cb9caef29b243;
    assign coff[676 ] = 64'h7ee34636ef29b243;
    assign coff[677 ] = 64'h4dd14c6e9a5f02f5;
    assign coff[678 ] = 64'hef29b243811cb9ca;
    assign coff[679 ] = 64'h9a5f02f5b22eb392;
    assign coff[680 ] = 64'h7bac1d31deff63f4;
    assign coff[681 ] = 64'h401d03219136d97d;
    assign coff[682 ] = 64'hdeff63f48453e2cf;
    assign coff[683 ] = 64'h9136d97dbfe2fcdf;
    assign coff[684 ] = 64'h6ec92683bfe2fcdf;
    assign coff[685 ] = 64'h21009c0c8453e2cf;
    assign coff[686 ] = 64'hbfe2fcdf9136d97d;
    assign coff[687 ] = 64'h8453e2cfdeff63f4;
    assign coff[688 ] = 64'h72db8828c7812572;
    assign coff[689 ] = 64'h2944a7a286d5c802;
    assign coff[690 ] = 64'hc78125728d2477d8;
    assign coff[691 ] = 64'h86d5c802d6bb585e;
    assign coff[692 ] = 64'h792a37fed6bb585e;
    assign coff[693 ] = 64'h387eda8e8d2477d8;
    assign coff[694 ] = 64'hd6bb585e86d5c802;
    assign coff[695 ] = 64'h8d2477d8c7812572;
    assign coff[696 ] = 64'h7fbc040af7c24f59;
    assign coff[697 ] = 64'h547ea0739fd9d22a;
    assign coff[698 ] = 64'hf7c24f598043fbf6;
    assign coff[699 ] = 64'h9fd9d22aab815f8d;
    assign coff[700 ] = 64'h60262dd6ab815f8d;
    assign coff[701 ] = 64'h083db0a78043fbf6;
    assign coff[702 ] = 64'hab815f8d9fd9d22a;
    assign coff[703 ] = 64'h8043fbf6f7c24f59;
    assign coff[704 ] = 64'h61b02876ad4a1aba;
    assign coff[705 ] = 64'h0a973ba580705b50;
    assign coff[706 ] = 64'had4a1aba9e4fd78a;
    assign coff[707 ] = 64'h80705b50f568c45b;
    assign coff[708 ] = 64'h7f8fa4b0f568c45b;
    assign coff[709 ] = 64'h52b5e5469e4fd78a;
    assign coff[710 ] = 64'hf568c45b80705b50;
    assign coff[711 ] = 64'h9e4fd78aad4a1aba;
    assign coff[712 ] = 64'h79e76ca7d8f81439;
    assign coff[713 ] = 64'h3a99a0578e33a9da;
    assign coff[714 ] = 64'hd8f8143986189359;
    assign coff[715 ] = 64'h8e33a9dac5665fa9;
    assign coff[716 ] = 64'h71cc5626c5665fa9;
    assign coff[717 ] = 64'h2707ebc786189359;
    assign coff[718 ] = 64'hc5665fa98e33a9da;
    assign coff[719 ] = 64'h86189359d8f81439;
    assign coff[720 ] = 64'h6ff27497c1efcdf3;
    assign coff[721 ] = 64'h2345eff884f4c2d4;
    assign coff[722 ] = 64'hc1efcdf3900d8b69;
    assign coff[723 ] = 64'h84f4c2d4dcba1008;
    assign coff[724 ] = 64'h7b0b3d2cdcba1008;
    assign coff[725 ] = 64'h3e10320d900d8b69;
    assign coff[726 ] = 64'hdcba100884f4c2d4;
    assign coff[727 ] = 64'h900d8b69c1efcdf3;
    assign coff[728 ] = 64'h7f2d1c0ef1805662;
    assign coff[729 ] = 64'h4faccfab9bd21af3;
    assign coff[730 ] = 64'hf180566280d2e3f2;
    assign coff[731 ] = 64'h9bd21af3b0533055;
    assign coff[732 ] = 64'h642de50db0533055;
    assign coff[733 ] = 64'h0e7fa99e80d2e3f2;
    assign coff[734 ] = 64'hb05330559bd21af3;
    assign coff[735 ] = 64'h80d2e3f2f1805662;
    assign coff[736 ] = 64'h69532442b7434a67;
    assign coff[737 ] = 64'h170afd8d82175990;
    assign coff[738 ] = 64'hb7434a6796acdbbe;
    assign coff[739 ] = 64'h82175990e8f50273;
    assign coff[740 ] = 64'h7de8a670e8f50273;
    assign coff[741 ] = 64'h48bcb59996acdbbe;
    assign coff[742 ] = 64'he8f5027382175990;
    assign coff[743 ] = 64'h96acdbbeb7434a67;
    assign coff[744 ] = 64'h7d24881be51b0e2a;
    assign coff[745 ] = 64'h4578db93947e5c33;
    assign coff[746 ] = 64'he51b0e2a82db77e5;
    assign coff[747 ] = 64'h947e5c33ba87246d;
    assign coff[748 ] = 64'h6b81a3cdba87246d;
    assign coff[749 ] = 64'h1ae4f1d682db77e5;
    assign coff[750 ] = 64'hba87246d947e5c33;
    assign coff[751 ] = 64'h82db77e5e51b0e2a;
    assign coff[752 ] = 64'h757dc5cacd355491;
    assign coff[753 ] = 64'h2f29ebcc890186f2;
    assign coff[754 ] = 64'hcd3554918a823a36;
    assign coff[755 ] = 64'h890186f2d0d61434;
    assign coff[756 ] = 64'h76fe790ed0d61434;
    assign coff[757 ] = 64'h32caab6f8a823a36;
    assign coff[758 ] = 64'hd0d61434890186f2;
    assign coff[759 ] = 64'h8a823a36cd355491;
    assign coff[760 ] = 64'h7ffc250ffe095d69;
    assign coff[761 ] = 64'h591c550ea41cd599;
    assign coff[762 ] = 64'hfe095d698003daf1;
    assign coff[763 ] = 64'ha41cd599a6e3aaf2;
    assign coff[764 ] = 64'h5be32a67a6e3aaf2;
    assign coff[765 ] = 64'h01f6a2978003daf1;
    assign coff[766 ] = 64'ha6e3aaf2a41cd599;
    assign coff[767 ] = 64'h8003daf1fe095d69;
    assign coff[768 ] = 64'h5c6eb258a7746ec0;
    assign coff[769 ] = 64'h02bfa9a480078e5e;
    assign coff[770 ] = 64'ha7746ec0a3914da8;
    assign coff[771 ] = 64'h80078e5efd40565c;
    assign coff[772 ] = 64'h7ff871a2fd40565c;
    assign coff[773 ] = 64'h588b9140a3914da8;
    assign coff[774 ] = 64'hfd40565c80078e5e;
    assign coff[775 ] = 64'ha3914da8a7746ec0;
    assign coff[776 ] = 64'h7747fbced191386e;
    assign coff[777 ] = 64'h3382fa888ad29394;
    assign coff[778 ] = 64'hd191386e88b80432;
    assign coff[779 ] = 64'h8ad29394cc7d0578;
    assign coff[780 ] = 64'h752d6c6ccc7d0578;
    assign coff[781 ] = 64'h2e6ec79288b80432;
    assign coff[782 ] = 64'hcc7d05788ad29394;
    assign coff[783 ] = 64'h88b80432d191386e;
    assign coff[784 ] = 64'h6bee3f62bb3058c0;
    assign coff[785 ] = 64'h1ba9633583065110;
    assign coff[786 ] = 64'hbb3058c09411c09e;
    assign coff[787 ] = 64'h83065110e4569ccb;
    assign coff[788 ] = 64'h7cf9aef0e4569ccb;
    assign coff[789 ] = 64'h44cfa7409411c09e;
    assign coff[790 ] = 64'he4569ccb83065110;
    assign coff[791 ] = 64'h9411c09ebb3058c0;
    assign coff[792 ] = 64'h7e0c3d29e9bae57d;
    assign coff[793 ] = 64'h4961cd33971f9ed7;
    assign coff[794 ] = 64'he9bae57d81f3c2d7;
    assign coff[795 ] = 64'h971f9ed7b69e32cd;
    assign coff[796 ] = 64'h68e06129b69e32cd;
    assign coff[797 ] = 64'h16451a8381f3c2d7;
    assign coff[798 ] = 64'hb69e32cd971f9ed7;
    assign coff[799 ] = 64'h81f3c2d7e9bae57d;
    assign coff[800 ] = 64'h64aa907fb0f0eeda;
    assign coff[801 ] = 64'h0f475bff80ea4712;
    assign coff[802 ] = 64'hb0f0eeda9b556f81;
    assign coff[803 ] = 64'h80ea4712f0b8a401;
    assign coff[804 ] = 64'h7f15b8eef0b8a401;
    assign coff[805 ] = 64'h4f0f11269b556f81;
    assign coff[806 ] = 64'hf0b8a40180ea4712;
    assign coff[807 ] = 64'h9b556f81b0f0eeda;
    assign coff[808 ] = 64'h7b420d7add7b8220;
    assign coff[809 ] = 64'h3ebfbdcd906f927c;
    assign coff[810 ] = 64'hdd7b822084bdf286;
    assign coff[811 ] = 64'h906f927cc1404233;
    assign coff[812 ] = 64'h6f906d84c1404233;
    assign coff[813 ] = 64'h22847de084bdf286;
    assign coff[814 ] = 64'hc1404233906f927c;
    assign coff[815 ] = 64'h84bdf286dd7b8220;
    assign coff[816 ] = 64'h7227d61cc61968a2;
    assign coff[817 ] = 64'h27c737d3865678eb;
    assign coff[818 ] = 64'hc61968a28dd829e4;
    assign coff[819 ] = 64'h865678ebd838c82d;
    assign coff[820 ] = 64'h79a98715d838c82d;
    assign coff[821 ] = 64'h39e6975e8dd829e4;
    assign coff[822 ] = 64'hd838c82d865678eb;
    assign coff[823 ] = 64'h8dd829e4c61968a2;
    assign coff[824 ] = 64'h7f9faa15f6313077;
    assign coff[825 ] = 64'h534ef1b59ed23bb9;
    assign coff[826 ] = 64'hf6313077806055eb;
    assign coff[827 ] = 64'h9ed23bb9acb10e4b;
    assign coff[828 ] = 64'h612dc447acb10e4b;
    assign coff[829 ] = 64'h09cecf89806055eb;
    assign coff[830 ] = 64'hacb10e4b9ed23bb9;
    assign coff[831 ] = 64'h806055ebf6313077;
    assign coff[832 ] = 64'h60aa7050ac18cf69;
    assign coff[833 ] = 64'h09064b3a80518b6b;
    assign coff[834 ] = 64'hac18cf699f558fb0;
    assign coff[835 ] = 64'h80518b6bf6f9b4c6;
    assign coff[836 ] = 64'h7fae7495f6f9b4c6;
    assign coff[837 ] = 64'h53e730979f558fb0;
    assign coff[838 ] = 64'hf6f9b4c680518b6b;
    assign coff[839 ] = 64'h9f558fb0ac18cf69;
    assign coff[840 ] = 64'h796a7554d779de47;
    assign coff[841 ] = 64'h3932ff878d7dc399;
    assign coff[842 ] = 64'hd779de4786958aac;
    assign coff[843 ] = 64'h8d7dc399c6cd0079;
    assign coff[844 ] = 64'h72823c67c6cd0079;
    assign coff[845 ] = 64'h288621b986958aac;
    assign coff[846 ] = 64'hc6cd00798d7dc399;
    assign coff[847 ] = 64'h86958aacd779de47;
    assign coff[848 ] = 64'h6f2d532cc0915148;
    assign coff[849 ] = 64'h21c2b69c84885258;
    assign coff[850 ] = 64'hc091514890d2acd4;
    assign coff[851 ] = 64'h84885258de3d4964;
    assign coff[852 ] = 64'h7b77ada8de3d4964;
    assign coff[853 ] = 64'h3f6eaeb890d2acd4;
    assign coff[854 ] = 64'hde3d496484885258;
    assign coff[855 ] = 64'h90d2acd4c0915148;
    assign coff[856 ] = 64'h7efd1c3ceff11753;
    assign coff[857 ] = 64'h4e708f8f9ad9bc71;
    assign coff[858 ] = 64'heff117538102e3c4;
    assign coff[859 ] = 64'h9ad9bc71b18f7071;
    assign coff[860 ] = 64'h6526438fb18f7071;
    assign coff[861 ] = 64'h100ee8ad8102e3c4;
    assign coff[862 ] = 64'hb18f70719ad9bc71;
    assign coff[863 ] = 64'h8102e3c4eff11753;
    assign coff[864 ] = 64'h686c9b4bb5f9d043;
    assign coff[865 ] = 64'h157f008681d16321;
    assign coff[866 ] = 64'hb5f9d043979364b5;
    assign coff[867 ] = 64'h81d16321ea80ff7a;
    assign coff[868 ] = 64'h7e2e9cdfea80ff7a;
    assign coff[869 ] = 64'h4a062fbd979364b5;
    assign coff[870 ] = 64'hea80ff7a81d16321;
    assign coff[871 ] = 64'h979364b5b5f9d043;
    assign coff[872 ] = 64'h7ccda169e3926fad;
    assign coff[873 ] = 64'h4425c92393a62f57;
    assign coff[874 ] = 64'he3926fad83325e97;
    assign coff[875 ] = 64'h93a62f57bbda36dd;
    assign coff[876 ] = 64'h6c59d0a9bbda36dd;
    assign coff[877 ] = 64'h1c6d905383325e97;
    assign coff[878 ] = 64'hbbda36dd93a62f57;
    assign coff[879 ] = 64'h83325e97e3926fad;
    assign coff[880 ] = 64'h74dbf1efcbc53579;
    assign coff[881 ] = 64'h2db330c7886fa7c2;
    assign coff[882 ] = 64'hcbc535798b240e11;
    assign coff[883 ] = 64'h886fa7c2d24ccf39;
    assign coff[884 ] = 64'h7790583ed24ccf39;
    assign coff[885 ] = 64'h343aca878b240e11;
    assign coff[886 ] = 64'hd24ccf39886fa7c2;
    assign coff[887 ] = 64'h8b240e11cbc53579;
    assign coff[888 ] = 64'h7ff38274fc775616;
    assign coff[889 ] = 64'h57f9f2f8a306a9c8;
    assign coff[890 ] = 64'hfc775616800c7d8c;
    assign coff[891 ] = 64'ha306a9c8a8060d08;
    assign coff[892 ] = 64'h5cf95638a8060d08;
    assign coff[893 ] = 64'h0388a9ea800c7d8c;
    assign coff[894 ] = 64'ha8060d08a306a9c8;
    assign coff[895 ] = 64'h800c7d8cfc775616;
    assign coff[896 ] = 64'h5e93dc1fa9bff8a8;
    assign coff[897 ] = 64'h05e36ea98022b114;
    assign coff[898 ] = 64'ha9bff8a8a16c23e1;
    assign coff[899 ] = 64'h8022b114fa1c9157;
    assign coff[900 ] = 64'h7fdd4eecfa1c9157;
    assign coff[901 ] = 64'h56400758a16c23e1;
    assign coff[902 ] = 64'hfa1c91578022b114;
    assign coff[903 ] = 64'ha16c23e1a9bff8a8;
    assign coff[904 ] = 64'h786280bfd48230e9;
    assign coff[905 ] = 64'h365f2e3b8c1f3c5d;
    assign coff[906 ] = 64'hd48230e9879d7f41;
    assign coff[907 ] = 64'h8c1f3c5dc9a0d1c5;
    assign coff[908 ] = 64'h73e0c3a3c9a0d1c5;
    assign coff[909 ] = 64'h2b7dcf17879d7f41;
    assign coff[910 ] = 64'hc9a0d1c58c1f3c5d;
    assign coff[911 ] = 64'h879d7f41d48230e9;
    assign coff[912 ] = 64'h6d963c54bddbbb7f;
    assign coff[913 ] = 64'h1eb86b4683bdbd0e;
    assign coff[914 ] = 64'hbddbbb7f9269c3ac;
    assign coff[915 ] = 64'h83bdbd0ee14794ba;
    assign coff[916 ] = 64'h7c4242f2e14794ba;
    assign coff[917 ] = 64'h422444819269c3ac;
    assign coff[918 ] = 64'he14794ba83bdbd0e;
    assign coff[919 ] = 64'h9269c3acbddbbb7f;
    assign coff[920 ] = 64'h7e8e6eb2ecd48407;
    assign coff[921 ] = 64'h4bef092d98f4bbbc;
    assign coff[922 ] = 64'hecd484078171914e;
    assign coff[923 ] = 64'h98f4bbbcb410f6d3;
    assign coff[924 ] = 64'h670b4444b410f6d3;
    assign coff[925 ] = 64'h132b7bf98171914e;
    assign coff[926 ] = 64'hb410f6d398f4bbbc;
    assign coff[927 ] = 64'h8171914eecd48407;
    assign coff[928 ] = 64'h66937e91b36f784f;
    assign coff[929 ] = 64'h1264994e815410d4;
    assign coff[930 ] = 64'hb36f784f996c816f;
    assign coff[931 ] = 64'h815410d4ed9b66b2;
    assign coff[932 ] = 64'h7eabef2ced9b66b2;
    assign coff[933 ] = 64'h4c9087b1996c816f;
    assign coff[934 ] = 64'hed9b66b2815410d4;
    assign coff[935 ] = 64'h996c816fb36f784f;
    assign coff[936 ] = 64'h7c116853e0848b7f;
    assign coff[937 ] = 64'h4177cfb1920265e4;
    assign coff[938 ] = 64'he0848b7f83ee97ad;
    assign coff[939 ] = 64'h920265e4be88304f;
    assign coff[940 ] = 64'h6dfd9a1cbe88304f;
    assign coff[941 ] = 64'h1f7b748183ee97ad;
    assign coff[942 ] = 64'hbe88304f920265e4;
    assign coff[943 ] = 64'h83ee97ade0848b7f;
    assign coff[944 ] = 64'h738acc9ec8eb0fd6;
    assign coff[945 ] = 64'h2ac080268759c2ef;
    assign coff[946 ] = 64'hc8eb0fd68c753362;
    assign coff[947 ] = 64'h8759c2efd53f7fda;
    assign coff[948 ] = 64'h78a63d11d53f7fda;
    assign coff[949 ] = 64'h3714f02a8c753362;
    assign coff[950 ] = 64'hd53f7fda8759c2ef;
    assign coff[951 ] = 64'h8c753362c8eb0fd6;
    assign coff[952 ] = 64'h7fd37153f953bf91;
    assign coff[953 ] = 64'h55ab0d46a0e51d8c;
    assign coff[954 ] = 64'hf953bf91802c8ead;
    assign coff[955 ] = 64'ha0e51d8caa54f2ba;
    assign coff[956 ] = 64'h5f1ae274aa54f2ba;
    assign coff[957 ] = 64'h06ac406f802c8ead;
    assign coff[958 ] = 64'haa54f2baa0e51d8c;
    assign coff[959 ] = 64'h802c8eadf953bf91;
    assign coff[960 ] = 64'h62b21c7bae7e965b;
    assign coff[961 ] = 64'h0c27c3898094162c;
    assign coff[962 ] = 64'hae7e965b9d4de385;
    assign coff[963 ] = 64'h8094162cf3d83c77;
    assign coff[964 ] = 64'h7f6be9d4f3d83c77;
    assign coff[965 ] = 64'h518169a59d4de385;
    assign coff[966 ] = 64'hf3d83c778094162c;
    assign coff[967 ] = 64'h9d4de385ae7e965b;
    assign coff[968 ] = 64'h7a5fb0d8da77cb63;
    assign coff[969 ] = 64'h3bfdfecd8eedf33b;
    assign coff[970 ] = 64'hda77cb6385a04f28;
    assign coff[971 ] = 64'h8eedf33bc4020133;
    assign coff[972 ] = 64'h71120cc5c4020133;
    assign coff[973 ] = 64'h2588349d85a04f28;
    assign coff[974 ] = 64'hc40201338eedf33b;
    assign coff[975 ] = 64'h85a04f28da77cb63;
    assign coff[976 ] = 64'h70b34525c350af26;
    assign coff[977 ] = 64'h24c7cd338565f1b0;
    assign coff[978 ] = 64'hc350af268f4cbadb;
    assign coff[979 ] = 64'h8565f1b0db3832cd;
    assign coff[980 ] = 64'h7a9a0e50db3832cd;
    assign coff[981 ] = 64'h3caf50da8f4cbadb;
    assign coff[982 ] = 64'hdb3832cd8565f1b0;
    assign coff[983 ] = 64'h8f4cbadbc350af26;
    assign coff[984 ] = 64'h7f5834b7f310248a;
    assign coff[985 ] = 64'h50e5fd6d9cce562c;
    assign coff[986 ] = 64'hf310248a80a7cb49;
    assign coff[987 ] = 64'h9cce562caf1a0293;
    assign coff[988 ] = 64'h6331a9d4af1a0293;
    assign coff[989 ] = 64'h0cefdb7680a7cb49;
    assign coff[990 ] = 64'haf1a02939cce562c;
    assign coff[991 ] = 64'h80a7cb49f310248a;
    assign coff[992 ] = 64'h6a359db9b88f926d;
    assign coff[993 ] = 64'h1896172882622aa6;
    assign coff[994 ] = 64'hb88f926d95ca6247;
    assign coff[995 ] = 64'h82622aa6e769e8d8;
    assign coff[996 ] = 64'h7d9dd55ae769e8d8;
    assign coff[997 ] = 64'h47706d9395ca6247;
    assign coff[998 ] = 64'he769e8d882622aa6;
    assign coff[999 ] = 64'h95ca6247b88f926d;
    assign coff[1000] = 64'h7d769bb5e6a4b616;
    assign coff[1001] = 64'h46c9405c955aae17;
    assign coff[1002] = 64'he6a4b6168289644b;
    assign coff[1003] = 64'h955aae17b936bfa4;
    assign coff[1004] = 64'h6aa551e9b936bfa4;
    assign coff[1005] = 64'h195b49ea8289644b;
    assign coff[1006] = 64'hb936bfa4955aae17;
    assign coff[1007] = 64'h8289644be6a4b616;
    assign coff[1008] = 64'h761b1211cea768f2;
    assign coff[1009] = 64'h309ed5568997fc8a;
    assign coff[1010] = 64'hcea768f289e4edef;
    assign coff[1011] = 64'h8997fc8acf612aaa;
    assign coff[1012] = 64'h76680376cf612aaa;
    assign coff[1013] = 64'h3158970e89e4edef;
    assign coff[1014] = 64'hcf612aaa8997fc8a;
    assign coff[1015] = 64'h89e4edefcea768f2;
    assign coff[1016] = 64'h7fffd886ff9b781d;
    assign coff[1017] = 64'h5a3b47aba5368c4b;
    assign coff[1018] = 64'hff9b781d8000277a;
    assign coff[1019] = 64'ha5368c4ba5c4b855;
    assign coff[1020] = 64'h5ac973b5a5c4b855;
    assign coff[1021] = 64'h006487e38000277a;
    assign coff[1022] = 64'ha5c4b855a5368c4b;
    assign coff[1023] = 64'h8000277aff9b781d;
    assign coff[1024] = 64'h5aecdbc5a5e8662f;
    assign coff[1025] = 64'h0096cbc1800058d4;
    assign coff[1026] = 64'ha5e8662fa513243b;
    assign coff[1027] = 64'h800058d4ff69343f;
    assign coff[1028] = 64'h7fffa72cff69343f;
    assign coff[1029] = 64'h5a1799d1a513243b;
    assign coff[1030] = 64'hff69343f800058d4;
    assign coff[1031] = 64'ha513243ba5e8662f;
    assign coff[1032] = 64'h767b1231cf8fade9;
    assign coff[1033] = 64'h3186f48789f857d8;
    assign coff[1034] = 64'hcf8fade98984edcf;
    assign coff[1035] = 64'h89f857d8ce790b79;
    assign coff[1036] = 64'h7607a828ce790b79;
    assign coff[1037] = 64'h307052178984edcf;
    assign coff[1038] = 64'hce790b7989f857d8;
    assign coff[1039] = 64'h8984edcfcf8fade9;
    assign coff[1040] = 64'h6ac115e2b960a64c;
    assign coff[1041] = 64'h198c8ce782936317;
    assign coff[1042] = 64'hb960a64c953eea1e;
    assign coff[1043] = 64'h82936317e6737319;
    assign coff[1044] = 64'h7d6c9ce9e6737319;
    assign coff[1045] = 64'h469f59b4953eea1e;
    assign coff[1046] = 64'he673731982936317;
    assign coff[1047] = 64'h953eea1eb960a64c;
    assign coff[1048] = 64'h7da77359e79b3f16;
    assign coff[1049] = 64'h479a1d6795e67850;
    assign coff[1050] = 64'he79b3f1682588ca7;
    assign coff[1051] = 64'h95e67850b865e299;
    assign coff[1052] = 64'h6a1987b0b865e299;
    assign coff[1053] = 64'h1864c0ea82588ca7;
    assign coff[1054] = 64'hb865e29995e67850;
    assign coff[1055] = 64'h82588ca7e79b3f16;
    assign coff[1056] = 64'h635166f9af40fce1;
    assign coff[1057] = 64'h0d21dc8780ace9ab;
    assign coff[1058] = 64'haf40fce19cae9907;
    assign coff[1059] = 64'h80ace9abf2de2379;
    assign coff[1060] = 64'h7f531655f2de2379;
    assign coff[1061] = 64'h50bf031f9cae9907;
    assign coff[1062] = 64'hf2de237980ace9ab;
    assign coff[1063] = 64'h9cae9907af40fce1;
    assign coff[1064] = 64'h7aa8766fdb685ae9;
    assign coff[1065] = 64'h3cdb8e098f649840;
    assign coff[1066] = 64'hdb685ae985578991;
    assign coff[1067] = 64'h8f649840c32471f7;
    assign coff[1068] = 64'h709b67c0c32471f7;
    assign coff[1069] = 64'h2497a51785578991;
    assign coff[1070] = 64'hc32471f78f649840;
    assign coff[1071] = 64'h85578991db685ae9;
    assign coff[1072] = 64'h7129931fc42e6ce8;
    assign coff[1073] = 64'h25b8401285af15b9;
    assign coff[1074] = 64'hc42e6ce88ed66ce1;
    assign coff[1075] = 64'h85af15b9da47bfee;
    assign coff[1076] = 64'h7a50ea47da47bfee;
    assign coff[1077] = 64'h3bd193188ed66ce1;
    assign coff[1078] = 64'hda47bfee85af15b9;
    assign coff[1079] = 64'h8ed66ce1c42e6ce8;
    assign coff[1080] = 64'h7f70a5fef40a4735;
    assign coff[1081] = 64'h51a825559d6decf4;
    assign coff[1082] = 64'hf40a4735808f5a02;
    assign coff[1083] = 64'h9d6decf4ae57daab;
    assign coff[1084] = 64'h6292130cae57daab;
    assign coff[1085] = 64'h0bf5b8cb808f5a02;
    assign coff[1086] = 64'hae57daab9d6decf4;
    assign coff[1087] = 64'h808f5a02f40a4735;
    assign coff[1088] = 64'h5f3c7f6baa7a5253;
    assign coff[1089] = 64'h06de7262802f375d;
    assign coff[1090] = 64'haa7a5253a0c38095;
    assign coff[1091] = 64'h802f375df9218d9e;
    assign coff[1092] = 64'h7fd0c8a3f9218d9e;
    assign coff[1093] = 64'h5585adada0c38095;
    assign coff[1094] = 64'hf9218d9e802f375d;
    assign coff[1095] = 64'ha0c38095aa7a5253;
    assign coff[1096] = 64'h78b6fda8d56ee424;
    assign coff[1097] = 64'h37424b7b8c8addb7;
    assign coff[1098] = 64'hd56ee42487490258;
    assign coff[1099] = 64'h8c8addb7c8bdb485;
    assign coff[1100] = 64'h73752249c8bdb485;
    assign coff[1101] = 64'h2a911bdc87490258;
    assign coff[1102] = 64'hc8bdb4858c8addb7;
    assign coff[1103] = 64'h87490258d56ee424;
    assign coff[1104] = 64'h6e174730beb366d1;
    assign coff[1105] = 64'h1fac2abf83fafe2e;
    assign coff[1106] = 64'hbeb366d191e8b8d0;
    assign coff[1107] = 64'h83fafe2ee053d541;
    assign coff[1108] = 64'h7c0501d2e053d541;
    assign coff[1109] = 64'h414c992f91e8b8d0;
    assign coff[1110] = 64'he053d54183fafe2e;
    assign coff[1111] = 64'h91e8b8d0beb366d1;
    assign coff[1112] = 64'h7eb31e78edcd2687;
    assign coff[1113] = 64'h4cb8c9dd998a9a74;
    assign coff[1114] = 64'hedcd2687814ce188;
    assign coff[1115] = 64'h998a9a74b3473623;
    assign coff[1116] = 64'h6675658cb3473623;
    assign coff[1117] = 64'h1232d979814ce188;
    assign coff[1118] = 64'hb3473623998a9a74;
    assign coff[1119] = 64'h814ce188edcd2687;
    assign coff[1120] = 64'h67290e02b43973ca;
    assign coff[1121] = 64'h135d2d538179223a;
    assign coff[1122] = 64'hb43973ca98d6f1fe;
    assign coff[1123] = 64'h8179223aeca2d2ad;
    assign coff[1124] = 64'h7e86ddc6eca2d2ad;
    assign coff[1125] = 64'h4bc68c3698d6f1fe;
    assign coff[1126] = 64'heca2d2ad8179223a;
    assign coff[1127] = 64'h98d6f1feb43973ca;
    assign coff[1128] = 64'h7c4e49b7e17862f3;
    assign coff[1129] = 64'h424f48459283c568;
    assign coff[1130] = 64'he17862f383b1b649;
    assign coff[1131] = 64'h9283c568bdb0b7bb;
    assign coff[1132] = 64'h6d7c3a98bdb0b7bb;
    assign coff[1133] = 64'h1e879d0d83b1b649;
    assign coff[1134] = 64'hbdb0b7bb9283c568;
    assign coff[1135] = 64'h83b1b649e17862f3;
    assign coff[1136] = 64'h73f614c0c9ce5748;
    assign coff[1137] = 64'h2bad122187ae9cc5;
    assign coff[1138] = 64'hc9ce57488c09eb40;
    assign coff[1139] = 64'h87ae9cc5d452eddf;
    assign coff[1140] = 64'h7851633bd452eddf;
    assign coff[1141] = 64'h3631a8b88c09eb40;
    assign coff[1142] = 64'hd452eddf87ae9cc5;
    assign coff[1143] = 64'h8c09eb40c9ce5748;
    assign coff[1144] = 64'h7fdf9508fa4ec821;
    assign coff[1145] = 64'h566524aaa18e09fa;
    assign coff[1146] = 64'hfa4ec82180206af8;
    assign coff[1147] = 64'ha18e09faa99adb56;
    assign coff[1148] = 64'h5e71f606a99adb56;
    assign coff[1149] = 64'h05b137df80206af8;
    assign coff[1150] = 64'ha99adb56a18e09fa;
    assign coff[1151] = 64'h80206af8fa4ec821;
    assign coff[1152] = 64'h5d1bdb65a82a9693;
    assign coff[1153] = 64'h03bae8b2800deaad;
    assign coff[1154] = 64'ha82a9693a2e4249b;
    assign coff[1155] = 64'h800deaadfc45174e;
    assign coff[1156] = 64'h7ff21553fc45174e;
    assign coff[1157] = 64'h57d5696da2e4249b;
    assign coff[1158] = 64'hfc45174e800deaad;
    assign coff[1159] = 64'ha2e4249ba82a9693;
    assign coff[1160] = 64'h77a24148d27bc69c;
    assign coff[1161] = 64'h3468aa768b3899c6;
    assign coff[1162] = 64'hd27bc69c885dbeb8;
    assign coff[1163] = 64'h8b3899c6cb97558a;
    assign coff[1164] = 64'h74c7663acb97558a;
    assign coff[1165] = 64'h2d843964885dbeb8;
    assign coff[1166] = 64'hcb97558a8b3899c6;
    assign coff[1167] = 64'h885dbeb8d27bc69c;
    assign coff[1168] = 64'h6c748b3fbc04c8ba;
    assign coff[1169] = 64'h1c9e90b8833d921b;
    assign coff[1170] = 64'hbc04c8ba938b74c1;
    assign coff[1171] = 64'h833d921be3616f48;
    assign coff[1172] = 64'h7cc26de5e3616f48;
    assign coff[1173] = 64'h43fb3746938b74c1;
    assign coff[1174] = 64'he3616f48833d921b;
    assign coff[1175] = 64'h938b74c1bc04c8ba;
    assign coff[1176] = 64'h7e37042aeab28e56;
    assign coff[1177] = 64'h4a2f2be697b07e7a;
    assign coff[1178] = 64'heab28e5681c8fbd6;
    assign coff[1179] = 64'h97b07e7ab5d0d41a;
    assign coff[1180] = 64'h684f8186b5d0d41a;
    assign coff[1181] = 64'h154d71aa81c8fbd6;
    assign coff[1182] = 64'hb5d0d41a97b07e7a;
    assign coff[1183] = 64'h81c8fbd6eab28e56;
    assign coff[1184] = 64'h6545095fb1b72f23;
    assign coff[1185] = 64'h1040c5bb81093be8;
    assign coff[1186] = 64'hb1b72f239abaf6a1;
    assign coff[1187] = 64'h81093be8efbf3a45;
    assign coff[1188] = 64'h7ef6c418efbf3a45;
    assign coff[1189] = 64'h4e48d0dd9abaf6a1;
    assign coff[1190] = 64'hefbf3a4581093be8;
    assign coff[1191] = 64'h9abaf6a1b1b72f23;
    assign coff[1192] = 64'h7b84e61fde6dc84b;
    assign coff[1193] = 64'h3f9a529090eb9e50;
    assign coff[1194] = 64'hde6dc84b847b19e1;
    assign coff[1195] = 64'h90eb9e50c065ad70;
    assign coff[1196] = 64'h6f1461b0c065ad70;
    assign coff[1197] = 64'h219237b5847b19e1;
    assign coff[1198] = 64'hc065ad7090eb9e50;
    assign coff[1199] = 64'h847b19e1de6dc84b;
    assign coff[1200] = 64'h7298a9ddc6f9fc8d;
    assign coff[1201] = 64'h28b5cca586a57df2;
    assign coff[1202] = 64'hc6f9fc8d8d675623;
    assign coff[1203] = 64'h86a57df2d74a335b;
    assign coff[1204] = 64'h795a820ed74a335b;
    assign coff[1205] = 64'h390603738d675623;
    assign coff[1206] = 64'hd74a335b86a57df2;
    assign coff[1207] = 64'h8d675623c6f9fc8d;
    assign coff[1208] = 64'h7fb1f5fcf72bd967;
    assign coff[1209] = 64'h540d20059f7689ff;
    assign coff[1210] = 64'hf72bd967804e0a04;
    assign coff[1211] = 64'h9f7689ffabf2dffb;
    assign coff[1212] = 64'h60897601abf2dffb;
    assign coff[1213] = 64'h08d42699804e0a04;
    assign coff[1214] = 64'habf2dffb9f7689ff;
    assign coff[1215] = 64'h804e0a04f72bd967;
    assign coff[1216] = 64'h614e73daacd73e30;
    assign coff[1217] = 64'h0a00ece8806439c0;
    assign coff[1218] = 64'hacd73e309eb18c26;
    assign coff[1219] = 64'h806439c0f5ff1318;
    assign coff[1220] = 64'h7f9bc640f5ff1318;
    assign coff[1221] = 64'h5328c1d09eb18c26;
    assign coff[1222] = 64'hf5ff1318806439c0;
    assign coff[1223] = 64'h9eb18c26acd73e30;
    assign coff[1224] = 64'h79b91ca4d868920f;
    assign coff[1225] = 64'h3a1367128deeef82;
    assign coff[1226] = 64'hd868920f8646e35c;
    assign coff[1227] = 64'h8deeef82c5ec98ee;
    assign coff[1228] = 64'h7211107ec5ec98ee;
    assign coff[1229] = 64'h27976df18646e35c;
    assign coff[1230] = 64'hc5ec98ee8deeef82;
    assign coff[1231] = 64'h8646e35cd868920f;
    assign coff[1232] = 64'h6fa90921c16c16b0;
    assign coff[1233] = 64'h22b4e27484cb8a1b;
    assign coff[1234] = 64'hc16c16b09056f6df;
    assign coff[1235] = 64'h84cb8a1bdd4b1d8c;
    assign coff[1236] = 64'h7b3475e5dd4b1d8c;
    assign coff[1237] = 64'h3e93e9509056f6df;
    assign coff[1238] = 64'hdd4b1d8c84cb8a1b;
    assign coff[1239] = 64'h9056f6dfc16c16b0;
    assign coff[1240] = 64'h7f1baf1ef0ea8d24;
    assign coff[1241] = 64'h4f3693209b748320;
    assign coff[1242] = 64'hf0ea8d2480e450e2;
    assign coff[1243] = 64'h9b748320b0c96ce0;
    assign coff[1244] = 64'h648b7ce0b0c96ce0;
    assign coff[1245] = 64'h0f1572dc80e450e2;
    assign coff[1246] = 64'hb0c96ce09b748320;
    assign coff[1247] = 64'h80e450e2f0ea8d24;
    assign coff[1248] = 64'h68fd2a3db6c767ca;
    assign coff[1249] = 64'h1676987f81fc8b60;
    assign coff[1250] = 64'hb6c767ca9702d5c3;
    assign coff[1251] = 64'h81fc8b60e9896781;
    assign coff[1252] = 64'h7e0374a0e9896781;
    assign coff[1253] = 64'h493898369702d5c3;
    assign coff[1254] = 64'he989678181fc8b60;
    assign coff[1255] = 64'h9702d5c3b6c767ca;
    assign coff[1256] = 64'h7d048228e487b2d0;
    assign coff[1257] = 64'h44fa0450942cce96;
    assign coff[1258] = 64'he487b2d082fb7dd8;
    assign coff[1259] = 64'h942cce96bb05fbb0;
    assign coff[1260] = 64'h6bd3316abb05fbb0;
    assign coff[1261] = 64'h1b784d3082fb7dd8;
    assign coff[1262] = 64'hbb05fbb0942cce96;
    assign coff[1263] = 64'h82fb7dd8e487b2d0;
    assign coff[1264] = 64'h75419de7ccab0d65;
    assign coff[1265] = 64'h2e9d9b7088ca4951;
    assign coff[1266] = 64'hccab0d658abe6219;
    assign coff[1267] = 64'h88ca4951d1626490;
    assign coff[1268] = 64'h7735b6afd1626490;
    assign coff[1269] = 64'h3354f29b8abe6219;
    assign coff[1270] = 64'hd162649088ca4951;
    assign coff[1271] = 64'h8abe6219ccab0d65;
    assign coff[1272] = 64'h7ff97c18fd729790;
    assign coff[1273] = 64'h58afd6bda3b41a50;
    assign coff[1274] = 64'hfd729790800683e8;
    assign coff[1275] = 64'ha3b41a50a7502943;
    assign coff[1276] = 64'h5c4be5b0a7502943;
    assign coff[1277] = 64'h028d6870800683e8;
    assign coff[1278] = 64'ha7502943a3b41a50;
    assign coff[1279] = 64'h800683e8fd729790;
    assign coff[1280] = 64'h5c0621b2a707c757;
    assign coff[1281] = 64'h0228e4e28004aa32;
    assign coff[1282] = 64'ha707c757a3f9de4e;
    assign coff[1283] = 64'h8004aa32fdd71b1e;
    assign coff[1284] = 64'h7ffb55cefdd71b1e;
    assign coff[1285] = 64'h58f838a9a3f9de4e;
    assign coff[1286] = 64'hfdd71b1e8004aa32;
    assign coff[1287] = 64'ha3f9de4ea707c757;
    assign coff[1288] = 64'h7710f54cd104d26b;
    assign coff[1289] = 64'h32f8cb078a963567;
    assign coff[1290] = 64'hd104d26b88ef0ab4;
    assign coff[1291] = 64'h8a963567cd0734f9;
    assign coff[1292] = 64'h7569ca99cd0734f9;
    assign coff[1293] = 64'h2efb2d9588ef0ab4;
    assign coff[1294] = 64'hcd0734f98a963567;
    assign coff[1295] = 64'h88ef0ab4d104d26b;
    assign coff[1296] = 64'h6b9ce39bbab16180;
    assign coff[1297] = 64'h1b16147982e61141;
    assign coff[1298] = 64'hbab1618094631c65;
    assign coff[1299] = 64'h82e61141e4e9eb87;
    assign coff[1300] = 64'h7d19eebfe4e9eb87;
    assign coff[1301] = 64'h454e9e8094631c65;
    assign coff[1302] = 64'he4e9eb8782e61141;
    assign coff[1303] = 64'h94631c65bab16180;
    assign coff[1304] = 64'h7df1a942e92675f4;
    assign coff[1305] = 64'h48e60c6296c97432;
    assign coff[1306] = 64'he92675f4820e56be;
    assign coff[1307] = 64'h96c97432b719f39e;
    assign coff[1308] = 64'h69368bceb719f39e;
    assign coff[1309] = 64'h16d98a0c820e56be;
    assign coff[1310] = 64'hb719f39e96c97432;
    assign coff[1311] = 64'h820e56bee92675f4;
    assign coff[1312] = 64'h644d2722b07a8d97;
    assign coff[1313] = 64'h0eb199a480d89f51;
    assign coff[1314] = 64'hb07a8d979bb2d8de;
    assign coff[1315] = 64'h80d89f51f14e665c;
    assign coff[1316] = 64'h7f2760aff14e665c;
    assign coff[1317] = 64'h4f8572699bb2d8de;
    assign coff[1318] = 64'hf14e665c80d89f51;
    assign coff[1319] = 64'h9bb2d8deb07a8d97;
    assign coff[1320] = 64'h7b190dbcdcea6478;
    assign coff[1321] = 64'h3e3c23699025f352;
    assign coff[1322] = 64'hdcea647884e6f244;
    assign coff[1323] = 64'h9025f352c1c3dc97;
    assign coff[1324] = 64'h6fda0caec1c3dc97;
    assign coff[1325] = 64'h23159b8884e6f244;
    assign coff[1326] = 64'hc1c3dc979025f352;
    assign coff[1327] = 64'h84e6f244dcea6478;
    assign coff[1328] = 64'h71e35080c593146a;
    assign coff[1329] = 64'h2737c7e38627f091;
    assign coff[1330] = 64'hc593146a8e1caf80;
    assign coff[1331] = 64'h8627f091d8c8381d;
    assign coff[1332] = 64'h79d80f6fd8c8381d;
    assign coff[1333] = 64'h3a6ceb968e1caf80;
    assign coff[1334] = 64'hd8c8381d8627f091;
    assign coff[1335] = 64'h8e1caf80c593146a;
    assign coff[1336] = 64'h7f93c38cf59add02;
    assign coff[1337] = 64'h52dc3b929e705a09;
    assign coff[1338] = 64'hf59add02806c3c74;
    assign coff[1339] = 64'h9e705a09ad23c46e;
    assign coff[1340] = 64'h618fa5f7ad23c46e;
    assign coff[1341] = 64'h0a6522fe806c3c74;
    assign coff[1342] = 64'had23c46e9e705a09;
    assign coff[1343] = 64'h806c3c74f59add02;
    assign coff[1344] = 64'h604754bfaba72807;
    assign coff[1345] = 64'h086fd94780474248;
    assign coff[1346] = 64'haba728079fb8ab41;
    assign coff[1347] = 64'h80474248f79026b9;
    assign coff[1348] = 64'h7fb8bdb8f79026b9;
    assign coff[1349] = 64'h5458d7f99fb8ab41;
    assign coff[1350] = 64'hf79026b980474248;
    assign coff[1351] = 64'h9fb8ab41aba72807;
    assign coff[1352] = 64'h793a6361d6eaf05f;
    assign coff[1353] = 64'h38abf0ef8d3ab03f;
    assign coff[1354] = 64'hd6eaf05f86c59c9f;
    assign coff[1355] = 64'h8d3ab03fc7540f11;
    assign coff[1356] = 64'h72c54fc1c7540f11;
    assign coff[1357] = 64'h29150fa186c59c9f;
    assign coff[1358] = 64'hc7540f118d3ab03f;
    assign coff[1359] = 64'h86c59c9fd6eaf05f;
    assign coff[1360] = 64'h6ee24b57c00e8336;
    assign coff[1361] = 64'h21312a658460e21a;
    assign coff[1362] = 64'hc00e8336911db4a9;
    assign coff[1363] = 64'h8460e21adeced59b;
    assign coff[1364] = 64'h7b9f1de6deced59b;
    assign coff[1365] = 64'h3ff17cca911db4a9;
    assign coff[1366] = 64'hdeced59b8460e21a;
    assign coff[1367] = 64'h911db4a9c00e8336;
    assign coff[1368] = 64'h7ee9d914ef5b87b5;
    assign coff[1369] = 64'h4df92f469a7d99de;
    assign coff[1370] = 64'hef5b87b5811626ec;
    assign coff[1371] = 64'h9a7d99deb206d0ba;
    assign coff[1372] = 64'h65826622b206d0ba;
    assign coff[1373] = 64'h10a4784b811626ec;
    assign coff[1374] = 64'hb206d0ba9a7d99de;
    assign coff[1375] = 64'h811626ecef5b87b5;
    assign coff[1376] = 64'h68151dbeb57efe22;
    assign coff[1377] = 64'h14ea4a1f81b867a5;
    assign coff[1378] = 64'hb57efe2297eae242;
    assign coff[1379] = 64'h81b867a5eb15b5e1;
    assign coff[1380] = 64'h7e47985beb15b5e1;
    assign coff[1381] = 64'h4a8101de97eae242;
    assign coff[1382] = 64'heb15b5e181b867a5;
    assign coff[1383] = 64'h97eae242b57efe22;
    assign coff[1384] = 64'h7cabcd28e2ff7bc3;
    assign coff[1385] = 64'h43a5f41e935631c5;
    assign coff[1386] = 64'he2ff7bc3835432d8;
    assign coff[1387] = 64'h935631c5bc5a0be2;
    assign coff[1388] = 64'h6ca9ce3bbc5a0be2;
    assign coff[1389] = 64'h1d00843d835432d8;
    assign coff[1390] = 64'hbc5a0be2935631c5;
    assign coff[1391] = 64'h835432d8e2ff7bc3;
    assign coff[1392] = 64'h749e18cdcb3badf3;
    assign coff[1393] = 64'h2d263596883a23ff;
    assign coff[1394] = 64'hcb3badf38b61e733;
    assign coff[1395] = 64'h883a23ffd2d9ca6a;
    assign coff[1396] = 64'h77c5dc01d2d9ca6a;
    assign coff[1397] = 64'h34c4520d8b61e733;
    assign coff[1398] = 64'hd2d9ca6a883a23ff;
    assign coff[1399] = 64'h8b61e733cb3badf3;
    assign coff[1400] = 64'h7feeffe1fbe09b80;
    assign coff[1401] = 64'h578c2dbaa29f4559;
    assign coff[1402] = 64'hfbe09b808011001f;
    assign coff[1403] = 64'ha29f4559a873d246;
    assign coff[1404] = 64'h5d60baa7a873d246;
    assign coff[1405] = 64'h041f64808011001f;
    assign coff[1406] = 64'ha873d246a29f4559;
    assign coff[1407] = 64'h8011001ffbe09b80;
    assign coff[1408] = 64'h5e2dfe29a950c8b0;
    assign coff[1409] = 64'h054cc7b1801c19ea;
    assign coff[1410] = 64'ha950c8b0a1d201d7;
    assign coff[1411] = 64'h801c19eafab3384f;
    assign coff[1412] = 64'h7fe3e616fab3384f;
    assign coff[1413] = 64'h56af3750a1d201d7;
    assign coff[1414] = 64'hfab3384f801c19ea;
    assign coff[1415] = 64'ha1d201d7a950c8b0;
    assign coff[1416] = 64'h782ef08bd3f47c06;
    assign coff[1417] = 64'h35d684a68bdf7eb0;
    assign coff[1418] = 64'hd3f47c0687d10f75;
    assign coff[1419] = 64'h8bdf7eb0ca297b5a;
    assign coff[1420] = 64'h74208150ca297b5a;
    assign coff[1421] = 64'h2c0b83fa87d10f75;
    assign coff[1422] = 64'hca297b5a8bdf7eb0;
    assign coff[1423] = 64'h87d10f75d3f47c06;
    assign coff[1424] = 64'h6d48047ebd5acee5;
    assign coff[1425] = 64'h1e25f2828399e244;
    assign coff[1426] = 64'hbd5acee592b7fb82;
    assign coff[1427] = 64'h8399e244e1da0d7e;
    assign coff[1428] = 64'h7c661dbce1da0d7e;
    assign coff[1429] = 64'h42a5311b92b7fb82;
    assign coff[1430] = 64'he1da0d7e8399e244;
    assign coff[1431] = 64'h92b7fb82bd5acee5;
    assign coff[1432] = 64'h7e778166ec3f78f6;
    assign coff[1433] = 64'h4b756f40989b8e40;
    assign coff[1434] = 64'hec3f78f681887e9a;
    assign coff[1435] = 64'h989b8e40b48a90c0;
    assign coff[1436] = 64'h676471c0b48a90c0;
    assign coff[1437] = 64'h13c0870a81887e9a;
    assign coff[1438] = 64'hb48a90c0989b8e40;
    assign coff[1439] = 64'h81887e9aec3f78f6;
    assign coff[1440] = 64'h66390422b2f6d550;
    assign coff[1441] = 64'h11cf516a813ebd90;
    assign coff[1442] = 64'hb2f6d55099c6fbde;
    assign coff[1443] = 64'h813ebd90ee30ae96;
    assign coff[1444] = 64'h7ec14270ee30ae96;
    assign coff[1445] = 64'h4d092ab099c6fbde;
    assign coff[1446] = 64'hee30ae96813ebd90;
    assign coff[1447] = 64'h99c6fbdeb2f6d550;
    assign coff[1448] = 64'h7bebfb70dff27773;
    assign coff[1449] = 64'h40f60dfb91b5919a;
    assign coff[1450] = 64'hdff2777384140490;
    assign coff[1451] = 64'h91b5919abf09f205;
    assign coff[1452] = 64'h6e4a6e66bf09f205;
    assign coff[1453] = 64'h200d888d84140490;
    assign coff[1454] = 64'hbf09f20591b5919a;
    assign coff[1455] = 64'h84140490dff27773;
    assign coff[1456] = 64'h73499838c863177b;
    assign coff[1457] = 64'h2a323f9e8727b905;
    assign coff[1458] = 64'hc863177b8cb667c8;
    assign coff[1459] = 64'h8727b905d5cdc062;
    assign coff[1460] = 64'h78d846fbd5cdc062;
    assign coff[1461] = 64'h379ce8858cb667c8;
    assign coff[1462] = 64'hd5cdc0628727b905;
    assign coff[1463] = 64'h8cb667c8c863177b;
    assign coff[1464] = 64'h7fcb3c23f8bd2cef;
    assign coff[1465] = 64'h553ac6eea08072ba;
    assign coff[1466] = 64'hf8bd2cef8034c3dd;
    assign coff[1467] = 64'ha08072baaac53912;
    assign coff[1468] = 64'h5f7f8d46aac53912;
    assign coff[1469] = 64'h0742d3118034c3dd;
    assign coff[1470] = 64'haac53912a08072ba;
    assign coff[1471] = 64'h8034c3ddf8bd2cef;
    assign coff[1472] = 64'h6251d298ae0a8916;
    assign coff[1473] = 64'h0b919dcf80861ca6;
    assign coff[1474] = 64'hae0a89169dae2d68;
    assign coff[1475] = 64'h80861ca6f46e6231;
    assign coff[1476] = 64'h7f79e35af46e6231;
    assign coff[1477] = 64'h51f576ea9dae2d68;
    assign coff[1478] = 64'hf46e623180861ca6;
    assign coff[1479] = 64'h9dae2d68ae0a8916;
    assign coff[1480] = 64'h7a332490d9e7ba7f;
    assign coff[1481] = 64'h3b78a0078ea7948c;
    assign coff[1482] = 64'hd9e7ba7f85ccdb70;
    assign coff[1483] = 64'h8ea7948cc4875ff9;
    assign coff[1484] = 64'h71586b74c4875ff9;
    assign coff[1485] = 64'h2618458185ccdb70;
    assign coff[1486] = 64'hc4875ff98ea7948c;
    assign coff[1487] = 64'h85ccdb70d9e7ba7f;
    assign coff[1488] = 64'h706b78e3c2cc13c7;
    assign coff[1489] = 64'h243743fa853af214;
    assign coff[1490] = 64'hc2cc13c78f94871d;
    assign coff[1491] = 64'h853af214dbc8bc06;
    assign coff[1492] = 64'h7ac50decdbc8bc06;
    assign coff[1493] = 64'h3d33ec398f94871d;
    assign coff[1494] = 64'hdbc8bc06853af214;
    assign coff[1495] = 64'h8f94871dc2cc13c7;
    assign coff[1496] = 64'h7f489eaaf27a2771;
    assign coff[1497] = 64'h5070e92f9c6f4cb6;
    assign coff[1498] = 64'hf27a277180b76156;
    assign coff[1499] = 64'h9c6f4cb6af8f16d1;
    assign coff[1500] = 64'h6390b34aaf8f16d1;
    assign coff[1501] = 64'h0d85d88f80b76156;
    assign coff[1502] = 64'haf8f16d19c6f4cb6;
    assign coff[1503] = 64'h80b76156f27a2771;
    assign coff[1504] = 64'h69e12a8cb812a41a;
    assign coff[1505] = 64'h1802092c82458acc;
    assign coff[1506] = 64'hb812a41a961ed574;
    assign coff[1507] = 64'h82458acce7fdf6d4;
    assign coff[1508] = 64'h7dba7534e7fdf6d4;
    assign coff[1509] = 64'h47ed5be6961ed574;
    assign coff[1510] = 64'he7fdf6d482458acc;
    assign coff[1511] = 64'h961ed574b812a41a;
    assign coff[1512] = 64'h7d58654de610f8f9;
    assign coff[1513] = 64'h464b6bbe95079394;
    assign coff[1514] = 64'he610f8f982a79ab3;
    assign coff[1515] = 64'h95079394b9b49442;
    assign coff[1516] = 64'h6af86c6cb9b49442;
    assign coff[1517] = 64'h19ef070782a79ab3;
    assign coff[1518] = 64'hb9b4944295079394;
    assign coff[1519] = 64'h82a79ab3e610f8f9;
    assign coff[1520] = 64'h75e09dbdce1c6777;
    assign coff[1521] = 64'h30133539895f072e;
    assign coff[1522] = 64'hce1c67778a1f6243;
    assign coff[1523] = 64'h895f072ecfeccac7;
    assign coff[1524] = 64'h76a0f8d2cfeccac7;
    assign coff[1525] = 64'h31e398898a1f6243;
    assign coff[1526] = 64'hcfeccac7895f072e;
    assign coff[1527] = 64'h8a1f6243ce1c6777;
    assign coff[1528] = 64'h7fff0943ff04acd0;
    assign coff[1529] = 64'h59d01475a4cc7e32;
    assign coff[1530] = 64'hff04acd08000f6bd;
    assign coff[1531] = 64'ha4cc7e32a62feb8b;
    assign coff[1532] = 64'h5b3381cea62feb8b;
    assign coff[1533] = 64'h00fb53308000f6bd;
    assign coff[1534] = 64'ha62feb8ba4cc7e32;
    assign coff[1535] = 64'h8000f6bdff04acd0;
    assign coff[1536] = 64'h5b79ef96a677a84e;
    assign coff[1537] = 64'h015fda038001e39b;
    assign coff[1538] = 64'ha677a84ea486106a;
    assign coff[1539] = 64'h8001e39bfea025fd;
    assign coff[1540] = 64'h7ffe1c65fea025fd;
    assign coff[1541] = 64'h598857b2a486106a;
    assign coff[1542] = 64'hfea025fd8001e39b;
    assign coff[1543] = 64'ha486106aa677a84e;
    assign coff[1544] = 64'h76c69647d04a054e;
    assign coff[1545] = 64'h32401dc68a46b564;
    assign coff[1546] = 64'hd04a054e893969b9;
    assign coff[1547] = 64'h8a46b564cdbfe23a;
    assign coff[1548] = 64'h75b94a9ccdbfe23a;
    assign coff[1549] = 64'h2fb5fab2893969b9;
    assign coff[1550] = 64'hcdbfe23a8a46b564;
    assign coff[1551] = 64'h893969b9d04a054e;
    assign coff[1552] = 64'h6b2f80fbba08ad95;
    assign coff[1553] = 64'h1a51712882bc1fa2;
    assign coff[1554] = 64'hba08ad9594d07f05;
    assign coff[1555] = 64'h82bc1fa2e5ae8ed8;
    assign coff[1556] = 64'h7d43e05ee5ae8ed8;
    assign coff[1557] = 64'h45f7526b94d07f05;
    assign coff[1558] = 64'he5ae8ed882bc1fa2;
    assign coff[1559] = 64'h94d07f05ba08ad95;
    assign coff[1560] = 64'h7dcd2981e860bd61;
    assign coff[1561] = 64'h48406e08965773e7;
    assign coff[1562] = 64'he860bd618232d67f;
    assign coff[1563] = 64'h965773e7b7bf91f8;
    assign coff[1564] = 64'h69a88c19b7bf91f8;
    assign coff[1565] = 64'h179f429f8232d67f;
    assign coff[1566] = 64'hb7bf91f8965773e7;
    assign coff[1567] = 64'h8232d67fe860bd61;
    assign coff[1568] = 64'h63cfc231afdd625f;
    assign coff[1569] = 64'h0de9cc4080c22784;
    assign coff[1570] = 64'hafdd625f9c303dcf;
    assign coff[1571] = 64'h80c22784f21633c0;
    assign coff[1572] = 64'h7f3dd87cf21633c0;
    assign coff[1573] = 64'h50229da19c303dcf;
    assign coff[1574] = 64'hf21633c080c22784;
    assign coff[1575] = 64'h9c303dcfafdd625f;
    assign coff[1576] = 64'h7ae159aedc293379;
    assign coff[1577] = 64'h3d8c24a88fc4bb53;
    assign coff[1578] = 64'hdc293379851ea652;
    assign coff[1579] = 64'h8fc4bb53c273db58;
    assign coff[1580] = 64'h703b44adc273db58;
    assign coff[1581] = 64'h23d6cc87851ea652;
    assign coff[1582] = 64'hc273db588fc4bb53;
    assign coff[1583] = 64'h851ea652dc293379;
    assign coff[1584] = 64'h7186fddec4e077b8;
    assign coff[1585] = 64'h2678337085eaec88;
    assign coff[1586] = 64'hc4e077b88e790222;
    assign coff[1587] = 64'h85eaec88d987cc90;
    assign coff[1588] = 64'h7a151378d987cc90;
    assign coff[1589] = 64'h3b1f88488e790222;
    assign coff[1590] = 64'hd987cc9085eaec88;
    assign coff[1591] = 64'h8e790222c4e077b8;
    assign coff[1592] = 64'h7f82d214f4d28451;
    assign coff[1593] = 64'h524295f09deeaa82;
    assign coff[1594] = 64'hf4d28451807d2dec;
    assign coff[1595] = 64'h9deeaa82adbd6a10;
    assign coff[1596] = 64'h6211557eadbd6a10;
    assign coff[1597] = 64'h0b2d7baf807d2dec;
    assign coff[1598] = 64'hadbd6a109deeaa82;
    assign coff[1599] = 64'h807d2decf4d28451;
    assign coff[1600] = 64'h5fc26038ab105464;
    assign coff[1601] = 64'h07a72f45803a9f31;
    assign coff[1602] = 64'hab105464a03d9fc8;
    assign coff[1603] = 64'h803a9f31f858d0bb;
    assign coff[1604] = 64'h7fc560cff858d0bb;
    assign coff[1605] = 64'h54efab9ca03d9fc8;
    assign coff[1606] = 64'hf858d0bb803a9f31;
    assign coff[1607] = 64'ha03d9fc8ab105464;
    assign coff[1608] = 64'h78f945c3d62cb6a8;
    assign coff[1609] = 64'h37f763418ce238f6;
    assign coff[1610] = 64'hd62cb6a88706ba3d;
    assign coff[1611] = 64'h8ce238f6c8089cbf;
    assign coff[1612] = 64'h731dc70ac8089cbf;
    assign coff[1613] = 64'h29d349588706ba3d;
    assign coff[1614] = 64'hc8089cbf8ce238f6;
    assign coff[1615] = 64'h8706ba3dd62cb6a8;
    assign coff[1616] = 64'h6e7d5193bf60a54a;
    assign coff[1617] = 64'h206ed295842d5762;
    assign coff[1618] = 64'hbf60a54a9182ae6d;
    assign coff[1619] = 64'h842d5762df912d6b;
    assign coff[1620] = 64'h7bd2a89edf912d6b;
    assign coff[1621] = 64'h409f5ab69182ae6d;
    assign coff[1622] = 64'hdf912d6b842d5762;
    assign coff[1623] = 64'h9182ae6dbf60a54a;
    assign coff[1624] = 64'h7ecf1837ee9441a0;
    assign coff[1625] = 64'h4d595bfe9a039c57;
    assign coff[1626] = 64'hee9441a08130e7c9;
    assign coff[1627] = 64'h9a039c57b2a6a402;
    assign coff[1628] = 64'h65fc63a9b2a6a402;
    assign coff[1629] = 64'h116bbe608130e7c9;
    assign coff[1630] = 64'hb2a6a4029a039c57;
    assign coff[1631] = 64'h8130e7c9ee9441a0;
    assign coff[1632] = 64'h679f95b7b4dbdc42;
    assign coff[1633] = 64'h1423d492819828fd;
    assign coff[1634] = 64'hb4dbdc4298606a49;
    assign coff[1635] = 64'h819828fdebdc2b6e;
    assign coff[1636] = 64'h7e67d703ebdc2b6e;
    assign coff[1637] = 64'h4b2423be98606a49;
    assign coff[1638] = 64'hebdc2b6e819828fd;
    assign coff[1639] = 64'h98606a49b4dbdc42;
    assign coff[1640] = 64'h7c7da505e23bcaa2;
    assign coff[1641] = 64'h42faf0d492ec7505;
    assign coff[1642] = 64'he23bcaa283825afb;
    assign coff[1643] = 64'h92ec7505bd050f2c;
    assign coff[1644] = 64'h6d138afbbd050f2c;
    assign coff[1645] = 64'h1dc4355e83825afb;
    assign coff[1646] = 64'hbd050f2c92ec7505;
    assign coff[1647] = 64'h83825afbe23bcaa2;
    assign coff[1648] = 64'h744aa63fca84c0a3;
    assign coff[1649] = 64'h2c69daa687f3cc48;
    assign coff[1650] = 64'hca84c0a38bb559c1;
    assign coff[1651] = 64'h87f3cc48d396255a;
    assign coff[1652] = 64'h780c33b8d396255a;
    assign coff[1653] = 64'h357b3f5d8bb559c1;
    assign coff[1654] = 64'hd396255a87f3cc48;
    assign coff[1655] = 64'h8bb559c1ca84c0a3;
    assign coff[1656] = 64'h7fe7e841fb17abc2;
    assign coff[1657] = 64'h56f9147ea21633cd;
    assign coff[1658] = 64'hfb17abc2801817bf;
    assign coff[1659] = 64'ha21633cda906eb82;
    assign coff[1660] = 64'h5de9cc33a906eb82;
    assign coff[1661] = 64'h04e8543e801817bf;
    assign coff[1662] = 64'ha906eb82a21633cd;
    assign coff[1663] = 64'h801817bffb17abc2;
    assign coff[1664] = 64'h5da5604fa8bd43fa;
    assign coff[1665] = 64'h0483ddc38014647b;
    assign coff[1666] = 64'ha8bd43faa25a9fb1;
    assign coff[1667] = 64'h8014647bfb7c223d;
    assign coff[1668] = 64'h7feb9b85fb7c223d;
    assign coff[1669] = 64'h5742bc06a25a9fb1;
    assign coff[1670] = 64'hfb7c223d8014647b;
    assign coff[1671] = 64'ha25a9fb1a8bd43fa;
    assign coff[1672] = 64'h77e92cd9d337ea12;
    assign coff[1673] = 64'h351fd9188b8b7c8f;
    assign coff[1674] = 64'hd337ea128816d327;
    assign coff[1675] = 64'h8b8b7c8fcae026e8;
    assign coff[1676] = 64'h74748371cae026e8;
    assign coff[1677] = 64'h2cc815ee8816d327;
    assign coff[1678] = 64'hcae026e88b8b7c8f;
    assign coff[1679] = 64'h8816d327d337ea12;
    assign coff[1680] = 64'h6cdece2fbcaf78c4;
    assign coff[1681] = 64'h1d6265dd836b207d;
    assign coff[1682] = 64'hbcaf78c4932131d1;
    assign coff[1683] = 64'h836b207de29d9a23;
    assign coff[1684] = 64'h7c94df83e29d9a23;
    assign coff[1685] = 64'h4350873c932131d1;
    assign coff[1686] = 64'he29d9a23836b207d;
    assign coff[1687] = 64'h932131d1bcaf78c4;
    assign coff[1688] = 64'h7e57dea7eb78ea52;
    assign coff[1689] = 64'h4ad2a9e29825863d;
    assign coff[1690] = 64'heb78ea5281a82159;
    assign coff[1691] = 64'h9825863db52d561e;
    assign coff[1692] = 64'h67da79c3b52d561e;
    assign coff[1693] = 64'h148715ae81a82159;
    assign coff[1694] = 64'hb52d561e9825863d;
    assign coff[1695] = 64'h81a82159eb78ea52;
    assign coff[1696] = 64'h65bf8447b256a26a;
    assign coff[1697] = 64'h110820968123603a;
    assign coff[1698] = 64'hb256a26a9a407bb9;
    assign coff[1699] = 64'h8123603aeef7df6a;
    assign coff[1700] = 64'h7edc9fc6eef7df6a;
    assign coff[1701] = 64'h4da95d969a407bb9;
    assign coff[1702] = 64'heef7df6a8123603a;
    assign coff[1703] = 64'h9a407bb9b256a26a;
    assign coff[1704] = 64'h7bb9096bdf2ff764;
    assign coff[1705] = 64'h40487f9491500f67;
    assign coff[1706] = 64'hdf2ff7648446f695;
    assign coff[1707] = 64'h91500f67bfb7806c;
    assign coff[1708] = 64'h6eaff099bfb7806c;
    assign coff[1709] = 64'h20d0089c8446f695;
    assign coff[1710] = 64'hbfb7806c91500f67;
    assign coff[1711] = 64'h8446f695df2ff764;
    assign coff[1712] = 64'h72f1aed9c7ae4489;
    assign coff[1713] = 64'h2974394686e60614;
    assign coff[1714] = 64'hc7ae44898d0e5127;
    assign coff[1715] = 64'h86e60614d68bc6ba;
    assign coff[1716] = 64'h7919f9ecd68bc6ba;
    assign coff[1717] = 64'h3851bb778d0e5127;
    assign coff[1718] = 64'hd68bc6ba86e60614;
    assign coff[1719] = 64'h8d0e5127c7ae4489;
    assign coff[1720] = 64'h7fbf36aaf7f4793e;
    assign coff[1721] = 64'h54a45be69ffb07e7;
    assign coff[1722] = 64'hf7f4793e8040c956;
    assign coff[1723] = 64'h9ffb07e7ab5ba41a;
    assign coff[1724] = 64'h6004f819ab5ba41a;
    assign coff[1725] = 64'h080b86c28040c956;
    assign coff[1726] = 64'hab5ba41a9ffb07e7;
    assign coff[1727] = 64'h8040c956f7f4793e;
    assign coff[1728] = 64'h61d09be5ad707dc8;
    assign coff[1729] = 64'h0ac952aa80748dd9;
    assign coff[1730] = 64'had707dc89e2f641b;
    assign coff[1731] = 64'h80748dd9f536ad56;
    assign coff[1732] = 64'h7f8b7227f536ad56;
    assign coff[1733] = 64'h528f82389e2f641b;
    assign coff[1734] = 64'hf536ad5680748dd9;
    assign coff[1735] = 64'h9e2f641bad707dc8;
    assign coff[1736] = 64'h79f6b711d927f65b;
    assign coff[1737] = 64'h3ac64c0f8e4ab5bf;
    assign coff[1738] = 64'hd927f65b860948ef;
    assign coff[1739] = 64'h8e4ab5bfc539b3f1;
    assign coff[1740] = 64'h71b54a41c539b3f1;
    assign coff[1741] = 64'h26d809a5860948ef;
    assign coff[1742] = 64'hc539b3f18e4ab5bf;
    assign coff[1743] = 64'h860948efd927f65b;
    assign coff[1744] = 64'h700acb3cc21bc8e1;
    assign coff[1745] = 64'h23763ef78502a65c;
    assign coff[1746] = 64'hc21bc8e18ff534c4;
    assign coff[1747] = 64'h8502a65cdc89c109;
    assign coff[1748] = 64'h7afd59a4dc89c109;
    assign coff[1749] = 64'h3de4371f8ff534c4;
    assign coff[1750] = 64'hdc89c1098502a65c;
    assign coff[1751] = 64'h8ff534c4c21bc8e1;
    assign coff[1752] = 64'h7f32c3d1f1b248a5;
    assign coff[1753] = 64'h4fd420a49bf16c7a;
    assign coff[1754] = 64'hf1b248a580cd3c2f;
    assign coff[1755] = 64'h9bf16c7ab02bdf5c;
    assign coff[1756] = 64'h640e9386b02bdf5c;
    assign coff[1757] = 64'h0e4db75b80cd3c2f;
    assign coff[1758] = 64'hb02bdf5c9bf16c7a;
    assign coff[1759] = 64'h80cd3c2ff1b248a5;
    assign coff[1760] = 64'h696fac78b76cac69;
    assign coff[1761] = 64'h173c6d8082206fcc;
    assign coff[1762] = 64'hb76cac6996905388;
    assign coff[1763] = 64'h82206fcce8c39280;
    assign coff[1764] = 64'h7ddf9034e8c39280;
    assign coff[1765] = 64'h4893539796905388;
    assign coff[1766] = 64'he8c3928082206fcc;
    assign coff[1767] = 64'h96905388b76cac69;
    assign coff[1768] = 64'h7d2f0e2be54c34f3;
    assign coff[1769] = 64'h45a30df09499ac95;
    assign coff[1770] = 64'he54c34f382d0f1d5;
    assign coff[1771] = 64'h9499ac95ba5cf210;
    assign coff[1772] = 64'h6b66536bba5cf210;
    assign coff[1773] = 64'h1ab3cb0d82d0f1d5;
    assign coff[1774] = 64'hba5cf2109499ac95;
    assign coff[1775] = 64'h82d0f1d5e54c34f3;
    assign coff[1776] = 64'h7591aeddcd637bfe;
    assign coff[1777] = 64'h2f58a2be89141589;
    assign coff[1778] = 64'hcd637bfe8a6e5123;
    assign coff[1779] = 64'h89141589d0a75d42;
    assign coff[1780] = 64'h76ebea77d0a75d42;
    assign coff[1781] = 64'h329c84028a6e5123;
    assign coff[1782] = 64'hd0a75d4289141589;
    assign coff[1783] = 64'h8a6e5123cd637bfe;
    assign coff[1784] = 64'h7ffce093fe3ba002;
    assign coff[1785] = 64'h594063b5a43fdb10;
    assign coff[1786] = 64'hfe3ba00280031f6d;
    assign coff[1787] = 64'ha43fdb10a6bf9c4b;
    assign coff[1788] = 64'h5bc024f0a6bf9c4b;
    assign coff[1789] = 64'h01c45ffe80031f6d;
    assign coff[1790] = 64'ha6bf9c4ba43fdb10;
    assign coff[1791] = 64'h80031f6dfe3ba002;
    assign coff[1792] = 64'h5c9170bfa798c1e5;
    assign coff[1793] = 64'h02f1ea6c8008ac90;
    assign coff[1794] = 64'ha798c1e5a36e8f41;
    assign coff[1795] = 64'h8008ac90fd0e1594;
    assign coff[1796] = 64'h7ff75370fd0e1594;
    assign coff[1797] = 64'h58673e1ba36e8f41;
    assign coff[1798] = 64'hfd0e15948008ac90;
    assign coff[1799] = 64'ha36e8f41a798c1e5;
    assign coff[1800] = 64'h775a2e89d1c01375;
    assign coff[1801] = 64'h33b0fa848ae6d720;
    assign coff[1802] = 64'hd1c0137588a5d177;
    assign coff[1803] = 64'h8ae6d720cc4f057c;
    assign coff[1804] = 64'h751928e0cc4f057c;
    assign coff[1805] = 64'h2e3fec8b88a5d177;
    assign coff[1806] = 64'hcc4f057c8ae6d720;
    assign coff[1807] = 64'h88a5d177d1c01375;
    assign coff[1808] = 64'h6c093cb6bb5ac06d;
    assign coff[1809] = 64'h1bda74f68311378d;
    assign coff[1810] = 64'hbb5ac06d93f6c34a;
    assign coff[1811] = 64'h8311378de4258b0a;
    assign coff[1812] = 64'h7ceec873e4258b0a;
    assign coff[1813] = 64'h44a53f9393f6c34a;
    assign coff[1814] = 64'he4258b0a8311378d;
    assign coff[1815] = 64'h93f6c34abb5ac06d;
    assign coff[1816] = 64'h7e14f242e9ec66e8;
    assign coff[1817] = 64'h498af6df973c7817;
    assign coff[1818] = 64'he9ec66e881eb0dbe;
    assign coff[1819] = 64'h973c7817b6750921;
    assign coff[1820] = 64'h68c387e9b6750921;
    assign coff[1821] = 64'h1613991881eb0dbe;
    assign coff[1822] = 64'hb6750921973c7817;
    assign coff[1823] = 64'h81eb0dbee9ec66e8;
    assign coff[1824] = 64'h64c99498b1187d05;
    assign coff[1825] = 64'h0f7942c780f050db;
    assign coff[1826] = 64'hb1187d059b366b68;
    assign coff[1827] = 64'h80f050dbf086bd39;
    assign coff[1828] = 64'h7f0faf25f086bd39;
    assign coff[1829] = 64'h4ee782fb9b366b68;
    assign coff[1830] = 64'hf086bd3980f050db;
    assign coff[1831] = 64'h9b366b68b1187d05;
    assign coff[1832] = 64'h7b4f920eddabec08;
    assign coff[1833] = 64'h3eeb889c90883f4d;
    assign coff[1834] = 64'hddabec0884b06df2;
    assign coff[1835] = 64'h90883f4dc1147764;
    assign coff[1836] = 64'h6f77c0b3c1147764;
    assign coff[1837] = 64'h225413f884b06df2;
    assign coff[1838] = 64'hc114776490883f4d;
    assign coff[1839] = 64'h84b06df2ddabec08;
    assign coff[1840] = 64'h723e8a20c6464144;
    assign coff[1841] = 64'h27f6fb928666213c;
    assign coff[1842] = 64'hc64641448dc175e0;
    assign coff[1843] = 64'h8666213cd809046e;
    assign coff[1844] = 64'h7999dec4d809046e;
    assign coff[1845] = 64'h39b9bebc8dc175e0;
    assign coff[1846] = 64'hd809046e8666213c;
    assign coff[1847] = 64'h8dc175e0c6464144;
    assign coff[1848] = 64'h7fa37a3cf6634f59;
    assign coff[1849] = 64'h537514c29ef2fa49;
    assign coff[1850] = 64'hf6634f59805c85c4;
    assign coff[1851] = 64'h9ef2fa49ac8aeb3e;
    assign coff[1852] = 64'h610d05b7ac8aeb3e;
    assign coff[1853] = 64'h099cb0a7805c85c4;
    assign coff[1854] = 64'hac8aeb3e9ef2fa49;
    assign coff[1855] = 64'h805c85c4f6634f59;
    assign coff[1856] = 64'h60cb5bb7ac3ecbc7;
    assign coff[1857] = 64'h09386e7880552084;
    assign coff[1858] = 64'hac3ecbc79f34a449;
    assign coff[1859] = 64'h80552084f6c79188;
    assign coff[1860] = 64'h7faadf7cf6c79188;
    assign coff[1861] = 64'h53c134399f34a449;
    assign coff[1862] = 64'hf6c7918880552084;
    assign coff[1863] = 64'h9f34a449ac3ecbc7;
    assign coff[1864] = 64'h797a55e0d7a98f73;
    assign coff[1865] = 64'h395ff2c98d9442b8;
    assign coff[1866] = 64'hd7a98f738685aa20;
    assign coff[1867] = 64'h8d9442b8c6a00d37;
    assign coff[1868] = 64'h726bbd48c6a00d37;
    assign coff[1869] = 64'h2856708d8685aa20;
    assign coff[1870] = 64'hc6a00d378d9442b8;
    assign coff[1871] = 64'h8685aa20d7a98f73;
    assign coff[1872] = 64'h6f463383c0bcfee7;
    assign coff[1873] = 64'h21f3304f84959dd9;
    assign coff[1874] = 64'hc0bcfee790b9cc7d;
    assign coff[1875] = 64'h84959dd9de0ccfb1;
    assign coff[1876] = 64'h7b6a6227de0ccfb1;
    assign coff[1877] = 64'h3f43011990b9cc7d;
    assign coff[1878] = 64'hde0ccfb184959dd9;
    assign coff[1879] = 64'h90b9cc7dc0bcfee7;
    assign coff[1880] = 64'h7f0360cbf022f6da;
    assign coff[1881] = 64'h4e9842299af891db;
    assign coff[1882] = 64'hf022f6da80fc9f35;
    assign coff[1883] = 64'h9af891dbb167bdd7;
    assign coff[1884] = 64'h65076e25b167bdd7;
    assign coff[1885] = 64'h0fdd092680fc9f35;
    assign coff[1886] = 64'hb167bdd79af891db;
    assign coff[1887] = 64'h80fc9f35f022f6da;
    assign coff[1888] = 64'h6889a4f6b622d7d6;
    assign coff[1889] = 64'h15b08c1281d9dde1;
    assign coff[1890] = 64'hb622d7d697765b0a;
    assign coff[1891] = 64'h81d9dde1ea4f73ee;
    assign coff[1892] = 64'h7e26221fea4f73ee;
    assign coff[1893] = 64'h49dd282a97765b0a;
    assign coff[1894] = 64'hea4f73ee81d9dde1;
    assign coff[1895] = 64'h97765b0ab622d7d6;
    assign coff[1896] = 64'h7cd8c1aee3c37474;
    assign coff[1897] = 64'h4450507e93c0faa3;
    assign coff[1898] = 64'he3c3747483273e52;
    assign coff[1899] = 64'h93c0faa3bbafaf82;
    assign coff[1900] = 64'h6c3f055dbbafaf82;
    assign coff[1901] = 64'h1c3c8b8c83273e52;
    assign coff[1902] = 64'hbbafaf8293c0faa3;
    assign coff[1903] = 64'h83273e52e3c37474;
    assign coff[1904] = 64'h74f06b9ecbf31d75;
    assign coff[1905] = 64'h2de2211e8881a33d;
    assign coff[1906] = 64'hcbf31d758b0f9462;
    assign coff[1907] = 64'h8881a33dd21ddee2;
    assign coff[1908] = 64'h777e5cc3d21ddee2;
    assign coff[1909] = 64'h340ce28b8b0f9462;
    assign coff[1910] = 64'hd21ddee28881a33d;
    assign coff[1911] = 64'h8b0f9462cbf31d75;
    assign coff[1912] = 64'h7ff4dbd9fca9956a;
    assign coff[1913] = 64'h581e6ef1a3293d4b;
    assign coff[1914] = 64'hfca9956a800b2427;
    assign coff[1915] = 64'ha3293d4ba7e1910f;
    assign coff[1916] = 64'h5cd6c2b5a7e1910f;
    assign coff[1917] = 64'h03566a96800b2427;
    assign coff[1918] = 64'ha7e1910fa3293d4b;
    assign coff[1919] = 64'h800b2427fca9956a;
    assign coff[1920] = 64'h5eb5b3a2a9e52347;
    assign coff[1921] = 64'h0615a48b80250ae7;
    assign coff[1922] = 64'ha9e52347a14a4c5e;
    assign coff[1923] = 64'h80250ae7f9ea5b75;
    assign coff[1924] = 64'h7fdaf519f9ea5b75;
    assign coff[1925] = 64'h561adcb9a14a4c5e;
    assign coff[1926] = 64'hf9ea5b7580250ae7;
    assign coff[1927] = 64'ha14a4c5ea9e52347;
    assign coff[1928] = 64'h78738bb3d4b17aa8;
    assign coff[1929] = 64'h368cab5c8c349f58;
    assign coff[1930] = 64'hd4b17aa8878c744d;
    assign coff[1931] = 64'h8c349f58c97354a4;
    assign coff[1932] = 64'h73cb60a8c97354a4;
    assign coff[1933] = 64'h2b4e8558878c744d;
    assign coff[1934] = 64'hc97354a48c349f58;
    assign coff[1935] = 64'h878c744dd4b17aa8;
    assign coff[1936] = 64'h6db02d29be06c977;
    assign coff[1937] = 64'h1ee934c383c9d6fc;
    assign coff[1938] = 64'hbe06c977924fd2d7;
    assign coff[1939] = 64'h83c9d6fce116cb3d;
    assign coff[1940] = 64'h7c362904e116cb3d;
    assign coff[1941] = 64'h41f93689924fd2d7;
    assign coff[1942] = 64'he116cb3d83c9d6fc;
    assign coff[1943] = 64'h924fd2d7be06c977;
    assign coff[1944] = 64'h7e95ec1aed063856;
    assign coff[1945] = 64'h4c177a6e9912955f;
    assign coff[1946] = 64'hed063856816a13e6;
    assign coff[1947] = 64'h9912955fb3e88592;
    assign coff[1948] = 64'h66ed6aa1b3e88592;
    assign coff[1949] = 64'h12f9c7aa816a13e6;
    assign coff[1950] = 64'hb3e885929912955f;
    assign coff[1951] = 64'h816a13e6ed063856;
    assign coff[1952] = 64'h66b187c3b397c649;
    assign coff[1953] = 64'h1296564d815b53a8;
    assign coff[1954] = 64'hb397c649994e783d;
    assign coff[1955] = 64'h815b53a8ed69a9b3;
    assign coff[1956] = 64'h7ea4ac58ed69a9b3;
    assign coff[1957] = 64'h4c6839b7994e783d;
    assign coff[1958] = 64'hed69a9b3815b53a8;
    assign coff[1959] = 64'h994e783db397c649;
    assign coff[1960] = 64'h7c1dbbb3e0b54698;
    assign coff[1961] = 64'h41a2fc1a921c23ef;
    assign coff[1962] = 64'he0b5469883e2444d;
    assign coff[1963] = 64'h921c23efbe5d03e6;
    assign coff[1964] = 64'h6de3dc11be5d03e6;
    assign coff[1965] = 64'h1f4ab96883e2444d;
    assign coff[1966] = 64'hbe5d03e6921c23ef;
    assign coff[1967] = 64'h83e2444de0b54698;
    assign coff[1968] = 64'h73a06522c91873a5;
    assign coff[1969] = 64'h2aefddd8876a9621;
    assign coff[1970] = 64'hc91873a58c5f9ade;
    assign coff[1971] = 64'h876a9621d5102228;
    assign coff[1972] = 64'h789569dfd5102228;
    assign coff[1973] = 64'h36e78c5b8c5f9ade;
    assign coff[1974] = 64'hd5102228876a9621;
    assign coff[1975] = 64'h8c5f9adec91873a5;
    assign coff[1976] = 64'h7fd6064cf985f28a;
    assign coff[1977] = 64'h55d05faaa106c92f;
    assign coff[1978] = 64'hf985f28a8029f9b4;
    assign coff[1979] = 64'ha106c92faa2fa056;
    assign coff[1980] = 64'h5ef936d1aa2fa056;
    assign coff[1981] = 64'h067a0d768029f9b4;
    assign coff[1982] = 64'haa2fa056a106c92f;
    assign coff[1983] = 64'h8029f9b4f985f28a;
    assign coff[1984] = 64'h62d216b3aea55e9e;
    assign coff[1985] = 64'h0c59cc688098e5fb;
    assign coff[1986] = 64'haea55e9e9d2de94d;
    assign coff[1987] = 64'h8098e5fbf3a63398;
    assign coff[1988] = 64'h7f671a05f3a63398;
    assign coff[1989] = 64'h515aa1629d2de94d;
    assign coff[1990] = 64'hf3a633988098e5fb;
    assign coff[1991] = 64'h9d2de94daea55e9e;
    assign coff[1992] = 64'h7a6e648adaa7dca1;
    assign coff[1993] = 64'h3c2a61428f058b04;
    assign coff[1994] = 64'hdaa7dca185919b76;
    assign coff[1995] = 64'h8f058b04c3d59ebe;
    assign coff[1996] = 64'h70fa74fcc3d59ebe;
    assign coff[1997] = 64'h2558235f85919b76;
    assign coff[1998] = 64'hc3d59ebe8f058b04;
    assign coff[1999] = 64'h85919b76daa7dca1;
    assign coff[2000] = 64'h70cb1128c37cf5b0;
    assign coff[2001] = 64'h24f7efa285746cb8;
    assign coff[2002] = 64'hc37cf5b08f34eed8;
    assign coff[2003] = 64'h85746cb8db08105e;
    assign coff[2004] = 64'h7a8b9348db08105e;
    assign coff[2005] = 64'h3c830a508f34eed8;
    assign coff[2006] = 64'hdb08105e85746cb8;
    assign coff[2007] = 64'h8f34eed8c37cf5b0;
    assign coff[2008] = 64'h7f5d3f75f342279b;
    assign coff[2009] = 64'h510ceb409cee229c;
    assign coff[2010] = 64'hf342279b80a2c08b;
    assign coff[2011] = 64'h9cee229caef314c0;
    assign coff[2012] = 64'h6311dd64aef314c0;
    assign coff[2013] = 64'h0cbdd86580a2c08b;
    assign coff[2014] = 64'haef314c09cee229c;
    assign coff[2015] = 64'h80a2c08bf342279b;
    assign coff[2016] = 64'h6a51a361b8b94d44;
    assign coff[2017] = 64'h18c7699b826bdc04;
    assign coff[2018] = 64'hb8b94d4495ae5c9f;
    assign coff[2019] = 64'h826bdc04e7389665;
    assign coff[2020] = 64'h7d9423fce7389665;
    assign coff[2021] = 64'h4746b2bc95ae5c9f;
    assign coff[2022] = 64'he7389665826bdc04;
    assign coff[2023] = 64'h95ae5c9fb8b94d44;
    assign coff[2024] = 64'h7d808728e6d5fcfc;
    assign coff[2025] = 64'h46f31c1a95768283;
    assign coff[2026] = 64'he6d5fcfc827f78d8;
    assign coff[2027] = 64'h95768283b90ce3e6;
    assign coff[2028] = 64'h6a897d7db90ce3e6;
    assign coff[2029] = 64'h192a0304827f78d8;
    assign coff[2030] = 64'hb90ce3e695768283;
    assign coff[2031] = 64'h827f78d8e6d5fcfc;
    assign coff[2032] = 64'h762e69c4ced5ce08;
    assign coff[2033] = 64'h30cd511589ab1d87;
    assign coff[2034] = 64'hced5ce0889d1963c;
    assign coff[2035] = 64'h89ab1d87cf32aeeb;
    assign coff[2036] = 64'h7654e279cf32aeeb;
    assign coff[2037] = 64'h312a31f889d1963c;
    assign coff[2038] = 64'hcf32aeeb89ab1d87;
    assign coff[2039] = 64'h89d1963cced5ce08;
    assign coff[2040] = 64'h7ffff621ffcdbc0b;
    assign coff[2041] = 64'h5a5ee79aa55a025b;
    assign coff[2042] = 64'hffcdbc0b800009df;
    assign coff[2043] = 64'ha55a025ba5a11866;
    assign coff[2044] = 64'h5aa5fda5a5a11866;
    assign coff[2045] = 64'h003243f5800009df;
    assign coff[2046] = 64'ha5a11866a55a025b;
    assign coff[2047] = 64'h800009dfffcdbc0b;
    assign coff[2048] = 64'h5ab7ba6ca5b2e6a0;
    assign coff[2049] = 64'h004b65ee80001635;
    assign coff[2050] = 64'ha5b2e6a0a5484594;
    assign coff[2051] = 64'h80001635ffb49a12;
    assign coff[2052] = 64'h7fffe9cbffb49a12;
    assign coff[2053] = 64'h5a4d1960a5484594;
    assign coff[2054] = 64'hffb49a1280001635;
    assign coff[2055] = 64'ha5484594a5b2e6a0;
    assign coff[2056] = 64'h765e7540cf49ebda;
    assign coff[2057] = 64'h3141657689db3fcf;
    assign coff[2058] = 64'hcf49ebda89a18ac0;
    assign coff[2059] = 64'h89db3fcfcebe9a8a;
    assign coff[2060] = 64'h7624c031cebe9a8a;
    assign coff[2061] = 64'h30b6142689a18ac0;
    assign coff[2062] = 64'hcebe9a8a89db3fcf;
    assign coff[2063] = 64'h89a18ac0cf49ebda;
    assign coff[2064] = 64'h6a9769c1b921d067;
    assign coff[2065] = 64'h1942a6f382846c26;
    assign coff[2066] = 64'hb921d0679568963f;
    assign coff[2067] = 64'h82846c26e6bd590d;
    assign coff[2068] = 64'h7d7b93dae6bd590d;
    assign coff[2069] = 64'h46de2f999568963f;
    assign coff[2070] = 64'he6bd590d82846c26;
    assign coff[2071] = 64'h9568963fb921d067;
    assign coff[2072] = 64'h7d98ff17e7513f25;
    assign coff[2073] = 64'h475b918895bc5d66;
    assign coff[2074] = 64'he7513f25826700e9;
    assign coff[2075] = 64'h95bc5d66b8a46e78;
    assign coff[2076] = 64'h6a43a29ab8a46e78;
    assign coff[2077] = 64'h18aec0db826700e9;
    assign coff[2078] = 64'hb8a46e7895bc5d66;
    assign coff[2079] = 64'h826700e9e7513f25;
    assign coff[2080] = 64'h6321c585af068a1a;
    assign coff[2081] = 64'h0cd6da2d80a54376;
    assign coff[2082] = 64'haf068a1a9cde3a7b;
    assign coff[2083] = 64'h80a54376f32925d3;
    assign coff[2084] = 64'h7f5abc8af32925d3;
    assign coff[2085] = 64'h50f975e69cde3a7b;
    assign coff[2086] = 64'hf32925d380a54376;
    assign coff[2087] = 64'h9cde3a7baf068a1a;
    assign coff[2088] = 64'h7a92d329db2020e0;
    assign coff[2089] = 64'h3c992ec08f40d2ad;
    assign coff[2090] = 64'hdb2020e0856d2cd7;
    assign coff[2091] = 64'h8f40d2adc366d140;
    assign coff[2092] = 64'h70bf2d53c366d140;
    assign coff[2093] = 64'h24dfdf20856d2cd7;
    assign coff[2094] = 64'hc366d1408f40d2ad;
    assign coff[2095] = 64'h856d2cd7db2020e0;
    assign coff[2096] = 64'h7106430ec3ebced0;
    assign coff[2097] = 64'h25702cb78598f2f3;
    assign coff[2098] = 64'hc3ebced08ef9bcf2;
    assign coff[2099] = 64'h8598f2f3da8fd349;
    assign coff[2100] = 64'h7a670d0dda8fd349;
    assign coff[2101] = 64'h3c1431308ef9bcf2;
    assign coff[2102] = 64'hda8fd3498598f2f3;
    assign coff[2103] = 64'h8ef9bcf2c3ebced0;
    assign coff[2104] = 64'h7f698461f3bf37cb;
    assign coff[2105] = 64'h516e07159d3de482;
    assign coff[2106] = 64'hf3bf37cb80967b9f;
    assign coff[2107] = 64'h9d3de482ae91f8eb;
    assign coff[2108] = 64'h62c21b7eae91f8eb;
    assign coff[2109] = 64'h0c40c83580967b9f;
    assign coff[2110] = 64'hae91f8eb9d3de482;
    assign coff[2111] = 64'h80967b9ff3bf37cb;
    assign coff[2112] = 64'h5f0a0e77aa4247e1;
    assign coff[2113] = 64'h06932713802b41ba;
    assign coff[2114] = 64'haa4247e1a0f5f189;
    assign coff[2115] = 64'h802b41baf96cd8ed;
    assign coff[2116] = 64'h7fd4be46f96cd8ed;
    assign coff[2117] = 64'h55bdb81fa0f5f189;
    assign coff[2118] = 64'hf96cd8ed802b41ba;
    assign coff[2119] = 64'ha0f5f189aa4247e1;
    assign coff[2120] = 64'h789dd5cbd527d02e;
    assign coff[2121] = 64'h36fe3f528c6a64e5;
    assign coff[2122] = 64'hd527d02e87622a35;
    assign coff[2123] = 64'h8c6a64e5c901c0ae;
    assign coff[2124] = 64'h73959b1bc901c0ae;
    assign coff[2125] = 64'h2ad82fd287622a35;
    assign coff[2126] = 64'hc901c0ae8c6a64e5;
    assign coff[2127] = 64'h87622a35d527d02e;
    assign coff[2128] = 64'h6df0bd35be7298d7;
    assign coff[2129] = 64'h1f63178f83e86b99;
    assign coff[2130] = 64'hbe7298d7920f42cb;
    assign coff[2131] = 64'h83e86b99e09ce871;
    assign coff[2132] = 64'h7c179467e09ce871;
    assign coff[2133] = 64'h418d6729920f42cb;
    assign coff[2134] = 64'he09ce87183e86b99;
    assign coff[2135] = 64'h920f42cbbe7298d7;
    assign coff[2136] = 64'h7ea85033ed8287d7;
    assign coff[2137] = 64'h4c7c622d995d7adc;
    assign coff[2138] = 64'hed8287d78157afcd;
    assign coff[2139] = 64'h995d7adcb3839dd3;
    assign coff[2140] = 64'h66a28524b3839dd3;
    assign coff[2141] = 64'h127d78298157afcd;
    assign coff[2142] = 64'hb3839dd3995d7adc;
    assign coff[2143] = 64'h8157afcded8287d7;
    assign coff[2144] = 64'h66fc596fb3fcbcbb;
    assign coff[2145] = 64'h1312a230816dd02a;
    assign coff[2146] = 64'hb3fcbcbb9903a691;
    assign coff[2147] = 64'h816dd02aeced5dd0;
    assign coff[2148] = 64'h7e922fd6eced5dd0;
    assign coff[2149] = 64'h4c0343459903a691;
    assign coff[2150] = 64'heced5dd0816dd02a;
    assign coff[2151] = 64'h9903a691b3fcbcbb;
    assign coff[2152] = 64'h7c3c3860e12f2f63;
    assign coff[2153] = 64'h420ebecb925cc924;
    assign coff[2154] = 64'he12f2f6383c3c7a0;
    assign coff[2155] = 64'h925cc924bdf14135;
    assign coff[2156] = 64'h6da336dcbdf14135;
    assign coff[2157] = 64'h1ed0d09d83c3c7a0;
    assign coff[2158] = 64'hbdf14135925cc924;
    assign coff[2159] = 64'h83c3c7a0e12f2f63;
    assign coff[2160] = 64'h73d61461c98a1227;
    assign coff[2161] = 64'h2b662b0e8794f774;
    assign coff[2162] = 64'hc98a12278c29eb9f;
    assign coff[2163] = 64'h8794f774d499d4f2;
    assign coff[2164] = 64'h786b088cd499d4f2;
    assign coff[2165] = 64'h3675edd98c29eb9f;
    assign coff[2166] = 64'hd499d4f28794f774;
    assign coff[2167] = 64'h8c29eb9fc98a1227;
    assign coff[2168] = 64'h7fdc247afa037648;
    assign coff[2169] = 64'h562d73b2a15b364d;
    assign coff[2170] = 64'hfa0376488023db86;
    assign coff[2171] = 64'ha15b364da9d28c4e;
    assign coff[2172] = 64'h5ea4c9b3a9d28c4e;
    assign coff[2173] = 64'h05fc89b88023db86;
    assign coff[2174] = 64'ha9d28c4ea15b364d;
    assign coff[2175] = 64'h8023db86fa037648;
    assign coff[2176] = 64'h5ce80e41a7f3cd59;
    assign coff[2177] = 64'h036f8a51800bce63;
    assign coff[2178] = 64'ha7f3cd59a317f1bf;
    assign coff[2179] = 64'h800bce63fc9075af;
    assign coff[2180] = 64'h7ff4319dfc9075af;
    assign coff[2181] = 64'h580c32a7a317f1bf;
    assign coff[2182] = 64'hfc9075af800bce63;
    assign coff[2183] = 64'ha317f1bfa7f3cd59;
    assign coff[2184] = 64'h77875cced235562b;
    assign coff[2185] = 64'h3423d78a8b19cef8;
    assign coff[2186] = 64'hd235562b8878a332;
    assign coff[2187] = 64'h8b19cef8cbdc2876;
    assign coff[2188] = 64'h74e63108cbdc2876;
    assign coff[2189] = 64'h2dcaa9d58878a332;
    assign coff[2190] = 64'hcbdc28768b19cef8;
    assign coff[2191] = 64'h8878a332d235562b;
    assign coff[2192] = 64'h6c4c6d1abbc4f1df;
    assign coff[2193] = 64'h1c550e7c832ccc0d;
    assign coff[2194] = 64'hbbc4f1df93b392e6;
    assign coff[2195] = 64'h832ccc0de3aaf184;
    assign coff[2196] = 64'h7cd333f3e3aaf184;
    assign coff[2197] = 64'h443b0e2193b392e6;
    assign coff[2198] = 64'he3aaf184832ccc0d;
    assign coff[2199] = 64'h93b392e6bbc4f1df;
    assign coff[2200] = 64'h7e2a61edea683949;
    assign coff[2201] = 64'h49f1ad619784dddc;
    assign coff[2202] = 64'hea68394981d59e13;
    assign coff[2203] = 64'h9784dddcb60e529f;
    assign coff[2204] = 64'h687b2224b60e529f;
    assign coff[2205] = 64'h1597c6b781d59e13;
    assign coff[2206] = 64'hb60e529f9784dddc;
    assign coff[2207] = 64'h81d59e13ea683949;
    assign coff[2208] = 64'h6516dacdb17b95a0;
    assign coff[2209] = 64'h0ff5f93880ffbf0a;
    assign coff[2210] = 64'hb17b95a09ae92533;
    assign coff[2211] = 64'h80ffbf0af00a06c8;
    assign coff[2212] = 64'h7f0040f6f00a06c8;
    assign coff[2213] = 64'h4e846a609ae92533;
    assign coff[2214] = 64'hf00a06c880ffbf0a;
    assign coff[2215] = 64'h9ae92533b17b95a0;
    assign coff[2216] = 64'h7b710a49de250be3;
    assign coff[2217] = 64'h3f58d92190c63a83;
    assign coff[2218] = 64'hde250be3848ef5b7;
    assign coff[2219] = 64'h90c63a83c0a726df;
    assign coff[2220] = 64'h6f39c57dc0a726df;
    assign coff[2221] = 64'h21daf41d848ef5b7;
    assign coff[2222] = 64'hc0a726df90c63a83;
    assign coff[2223] = 64'h848ef5b7de250be3;
    assign coff[2224] = 64'h7276ff0dc6b685bd;
    assign coff[2225] = 64'h286e49ea868d980e;
    assign coff[2226] = 64'hc6b685bd8d8900f3;
    assign coff[2227] = 64'h868d980ed791b616;
    assign coff[2228] = 64'h797267f2d791b616;
    assign coff[2229] = 64'h39497a438d8900f3;
    assign coff[2230] = 64'hd791b616868d980e;
    assign coff[2231] = 64'h8d8900f3c6b685bd;
    assign coff[2232] = 64'h7facac7ff6e0a2fa;
    assign coff[2233] = 64'h53d434069f45181f;
    assign coff[2234] = 64'hf6e0a2fa80535381;
    assign coff[2235] = 64'h9f45181fac2bcbfa;
    assign coff[2236] = 64'h60bae7e1ac2bcbfa;
    assign coff[2237] = 64'h091f5d0680535381;
    assign coff[2238] = 64'hac2bcbfa9f45181f;
    assign coff[2239] = 64'h80535381f6e0a2fa;
    assign coff[2240] = 64'h611d66deac9dfb29;
    assign coff[2241] = 64'h09b5c048805e6b62;
    assign coff[2242] = 64'hac9dfb299ee29922;
    assign coff[2243] = 64'h805e6b62f64a3fb8;
    assign coff[2244] = 64'h7fa1949ef64a3fb8;
    assign coff[2245] = 64'h536204d79ee29922;
    assign coff[2246] = 64'hf64a3fb8805e6b62;
    assign coff[2247] = 64'h9ee29922ac9dfb29;
    assign coff[2248] = 64'h79a1b545d820e589;
    assign coff[2249] = 64'h39d02c2a8dcccdaf;
    assign coff[2250] = 64'hd820e589865e4abb;
    assign coff[2251] = 64'h8dcccdafc62fd3d6;
    assign coff[2252] = 64'h72333251c62fd3d6;
    assign coff[2253] = 64'h27df1a77865e4abb;
    assign coff[2254] = 64'hc62fd3d68dcccdaf;
    assign coff[2255] = 64'h865e4abbd820e589;
    assign coff[2256] = 64'h6f841942c12a5b95;
    assign coff[2257] = 64'h226c499684b72ddb;
    assign coff[2258] = 64'hc12a5b95907be6be;
    assign coff[2259] = 64'h84b72ddbdd93b66a;
    assign coff[2260] = 64'h7b48d225dd93b66a;
    assign coff[2261] = 64'h3ed5a46b907be6be;
    assign coff[2262] = 64'hdd93b66a84b72ddb;
    assign coff[2263] = 64'h907be6bec12a5b95;
    assign coff[2264] = 64'h7f12b67cf09fb051;
    assign coff[2265] = 64'h4efb4b969b45eb83;
    assign coff[2266] = 64'hf09fb05180ed4984;
    assign coff[2267] = 64'h9b45eb83b104b46a;
    assign coff[2268] = 64'h64ba147db104b46a;
    assign coff[2269] = 64'h0f604faf80ed4984;
    assign coff[2270] = 64'hb104b46a9b45eb83;
    assign coff[2271] = 64'h80ed4984f09fb051;
    assign coff[2272] = 64'h68d1f68fb6899c8d;
    assign coff[2273] = 64'h162c5a3b81ef65dc;
    assign coff[2274] = 64'hb6899c8d972e0971;
    assign coff[2275] = 64'h81ef65dce9d3a5c5;
    assign coff[2276] = 64'h7e109a24e9d3a5c5;
    assign coff[2277] = 64'h49766373972e0971;
    assign coff[2278] = 64'he9d3a5c581ef65dc;
    assign coff[2279] = 64'h972e0971b6899c8d;
    assign coff[2280] = 64'h7cf43e1ae43e1362;
    assign coff[2281] = 64'h44ba74bd94043fdf;
    assign coff[2282] = 64'he43e1362830bc1e6;
    assign coff[2283] = 64'h94043fdfbb458b43;
    assign coff[2284] = 64'h6bfbc021bb458b43;
    assign coff[2285] = 64'h1bc1ec9e830bc1e6;
    assign coff[2286] = 64'hbb458b4394043fdf;
    assign coff[2287] = 64'h830bc1e6e43e1362;
    assign coff[2288] = 64'h75234ce8cc66047b;
    assign coff[2289] = 64'h2e575af388aee888;
    assign coff[2290] = 64'hcc66047b8adcb318;
    assign coff[2291] = 64'h88aee888d1a8a50d;
    assign coff[2292] = 64'h77511778d1a8a50d;
    assign coff[2293] = 64'h3399fb858adcb318;
    assign coff[2294] = 64'hd1a8a50d88aee888;
    assign coff[2295] = 64'h8adcb318cc66047b;
    assign coff[2296] = 64'h7ff7e500fd2735ea;
    assign coff[2297] = 64'h58796962a37fecac;
    assign coff[2298] = 64'hfd2735ea80081b00;
    assign coff[2299] = 64'ha37fecaca786969e;
    assign coff[2300] = 64'h5c801354a786969e;
    assign coff[2301] = 64'h02d8ca1680081b00;
    assign coff[2302] = 64'ha786969ea37fecac;
    assign coff[2303] = 64'h80081b00fd2735ea;
    assign coff[2304] = 64'h5bd1a971a6d1a1e7;
    assign coff[2305] = 64'h01dd815480037ab7;
    assign coff[2306] = 64'ha6d1a1e7a42e568f;
    assign coff[2307] = 64'h80037ab7fe227eac;
    assign coff[2308] = 64'h7ffc8549fe227eac;
    assign coff[2309] = 64'h592e5e19a42e568f;
    assign coff[2310] = 64'hfe227eac80037ab7;
    assign coff[2311] = 64'ha42e568fa6d1a1e7;
    assign coff[2312] = 64'h76f5340ed0beb7d2;
    assign coff[2313] = 64'h32b398b38a784368;
    assign coff[2314] = 64'hd0beb7d2890acbf2;
    assign coff[2315] = 64'h8a784368cd4c674d;
    assign coff[2316] = 64'h7587bc98cd4c674d;
    assign coff[2317] = 64'h2f41482e890acbf2;
    assign coff[2318] = 64'hcd4c674d8a784368;
    assign coff[2319] = 64'h890acbf2d0beb7d2;
    assign coff[2320] = 64'h6b73fdaeba7209e7;
    assign coff[2321] = 64'h1acc5ef682d63274;
    assign coff[2322] = 64'hba7209e7948c0252;
    assign coff[2323] = 64'h82d63274e533a10a;
    assign coff[2324] = 64'h7d29cd8ce533a10a;
    assign coff[2325] = 64'h458df619948c0252;
    assign coff[2326] = 64'he533a10a82d63274;
    assign coff[2327] = 64'h948c0252ba7209e7;
    assign coff[2328] = 64'h7de41dc0e8dc4a07;
    assign coff[2329] = 64'h48a805ff969e959b;
    assign coff[2330] = 64'he8dc4a07821be240;
    assign coff[2331] = 64'h969e959bb757fa01;
    assign coff[2332] = 64'h69616a65b757fa01;
    assign coff[2333] = 64'h1723b5f9821be240;
    assign coff[2334] = 64'hb757fa01969e959b;
    assign coff[2335] = 64'h821be240e8dc4a07;
    assign coff[2336] = 64'h641e3e38b03f864f;
    assign coff[2337] = 64'h0e66b0c380d00d9d;
    assign coff[2338] = 64'hb03f864f9be1c1c8;
    assign coff[2339] = 64'h80d00d9df1994f3d;
    assign coff[2340] = 64'h7f2ff263f1994f3d;
    assign coff[2341] = 64'h4fc079b19be1c1c8;
    assign coff[2342] = 64'hf1994f3d80d00d9d;
    assign coff[2343] = 64'h9be1c1c8b03f864f;
    assign coff[2344] = 64'h7b044dc7dca1e7da;
    assign coff[2345] = 64'h3dfa35c890015dee;
    assign coff[2346] = 64'hdca1e7da84fbb239;
    assign coff[2347] = 64'h90015deec205ca38;
    assign coff[2348] = 64'h6ffea212c205ca38;
    assign coff[2349] = 64'h235e182684fbb239;
    assign coff[2350] = 64'hc205ca3890015dee;
    assign coff[2351] = 64'h84fbb239dca1e7da;
    assign coff[2352] = 64'h71c0d265c55008ab;
    assign coff[2353] = 64'h26effb768610ebca;
    assign coff[2354] = 64'hc55008ab8e3f2d9b;
    assign coff[2355] = 64'h8610ebcad910048a;
    assign coff[2356] = 64'h79ef1436d910048a;
    assign coff[2357] = 64'h3aaff7558e3f2d9b;
    assign coff[2358] = 64'hd910048a8610ebca;
    assign coff[2359] = 64'h8e3f2d9bc55008ab;
    assign coff[2360] = 64'h7f8d8de1f54fb8a4;
    assign coff[2361] = 64'h52a2b5569e3f9bf0;
    assign coff[2362] = 64'hf54fb8a48072721f;
    assign coff[2363] = 64'h9e3f9bf0ad5d4aaa;
    assign coff[2364] = 64'h61c06410ad5d4aaa;
    assign coff[2365] = 64'h0ab0475c8072721f;
    assign coff[2366] = 64'had5d4aaa9e3f9bf0;
    assign coff[2367] = 64'h8072721ff54fb8a4;
    assign coff[2368] = 64'h601594d1ab6e8032;
    assign coff[2369] = 64'h08249bdd80426030;
    assign coff[2370] = 64'hab6e80329fea6b2f;
    assign coff[2371] = 64'h80426030f7db6423;
    assign coff[2372] = 64'h7fbd9fd0f7db6423;
    assign coff[2373] = 64'h54917fce9fea6b2f;
    assign coff[2374] = 64'hf7db642380426030;
    assign coff[2375] = 64'h9fea6b2fab6e8032;
    assign coff[2376] = 64'h79221b4bd6a38ec0;
    assign coff[2377] = 64'h38684c198d196249;
    assign coff[2378] = 64'hd6a38ec086dde4b5;
    assign coff[2379] = 64'h8d196249c797b3e7;
    assign coff[2380] = 64'h72e69db7c797b3e7;
    assign coff[2381] = 64'h295c714086dde4b5;
    assign coff[2382] = 64'hc797b3e78d196249;
    assign coff[2383] = 64'h86dde4b5d6a38ec0;
    assign coff[2384] = 64'h6ebc8db0bfcd3d69;
    assign coff[2385] = 64'h20e852f6844d6a50;
    assign coff[2386] = 64'hbfcd3d6991437250;
    assign coff[2387] = 64'h844d6a50df17ad0a;
    assign coff[2388] = 64'h7bb295b0df17ad0a;
    assign coff[2389] = 64'h4032c29791437250;
    assign coff[2390] = 64'hdf17ad0a844d6a50;
    assign coff[2391] = 64'h91437250bfcd3d69;
    assign coff[2392] = 64'h7edff570ef10c883;
    assign coff[2393] = 64'h4dbd56829a4fbd61;
    assign coff[2394] = 64'hef10c88381200a90;
    assign coff[2395] = 64'h9a4fbd61b242a97e;
    assign coff[2396] = 64'h65b0429fb242a97e;
    assign coff[2397] = 64'h10ef377d81200a90;
    assign coff[2398] = 64'hb242a97e9a4fbd61;
    assign coff[2399] = 64'h81200a90ef10c883;
    assign coff[2400] = 64'h67e928c5b541bbcd;
    assign coff[2401] = 64'h149fe3fc81ac2b9e;
    assign coff[2402] = 64'hb541bbcd9816d73b;
    assign coff[2403] = 64'h81ac2b9eeb601c04;
    assign coff[2404] = 64'h7e53d462eb601c04;
    assign coff[2405] = 64'h4abe44339816d73b;
    assign coff[2406] = 64'heb601c0481ac2b9e;
    assign coff[2407] = 64'h9816d73bb541bbcd;
    assign coff[2408] = 64'h7c9aa221e2b610da;
    assign coff[2409] = 64'h4365e65b932e6b84;
    assign coff[2410] = 64'he2b610da83655ddf;
    assign coff[2411] = 64'h932e6b84bc9a19a5;
    assign coff[2412] = 64'h6cd1947cbc9a19a5;
    assign coff[2413] = 64'h1d49ef2683655ddf;
    assign coff[2414] = 64'hbc9a19a5932e6b84;
    assign coff[2415] = 64'h83655ddfe2b610da;
    assign coff[2416] = 64'h747eef85caf7059a;
    assign coff[2417] = 64'h2cdfa071881fa06f;
    assign coff[2418] = 64'hcaf7059a8b81107b;
    assign coff[2419] = 64'h881fa06fd3205f8f;
    assign coff[2420] = 64'h77e05f91d3205f8f;
    assign coff[2421] = 64'h3508fa668b81107b;
    assign coff[2422] = 64'hd3205f8f881fa06f;
    assign coff[2423] = 64'h8b81107bcaf7059a;
    assign coff[2424] = 64'h7fec7c02fb95404d;
    assign coff[2425] = 64'h57551d80a26bc3b2;
    assign coff[2426] = 64'hfb95404d801383fe;
    assign coff[2427] = 64'ha26bc3b2a8aae280;
    assign coff[2428] = 64'h5d943c4ea8aae280;
    assign coff[2429] = 64'h046abfb3801383fe;
    assign coff[2430] = 64'ha8aae280a26bc3b2;
    assign coff[2431] = 64'h801383fefb95404d;
    assign coff[2432] = 64'h5dfade20a9195dc7;
    assign coff[2433] = 64'h05017165801910e4;
    assign coff[2434] = 64'ha9195dc7a20521e0;
    assign coff[2435] = 64'h801910e4fafe8e9b;
    assign coff[2436] = 64'h7fe6ef1cfafe8e9b;
    assign coff[2437] = 64'h56e6a239a20521e0;
    assign coff[2438] = 64'hfafe8e9b801910e4;
    assign coff[2439] = 64'ha20521e0a9195dc7;
    assign coff[2440] = 64'h7814e9dfd3adb876;
    assign coff[2441] = 64'h359213c98bbfdc44;
    assign coff[2442] = 64'hd3adb87687eb1621;
    assign coff[2443] = 64'h8bbfdc44ca6dec37;
    assign coff[2444] = 64'h744023bcca6dec37;
    assign coff[2445] = 64'h2c52478a87eb1621;
    assign coff[2446] = 64'hca6dec378bbfdc44;
    assign coff[2447] = 64'h87eb1621d3adb876;
    assign coff[2448] = 64'h6d20afacbd1a7b3d;
    assign coff[2449] = 64'h1ddca6628388359b;
    assign coff[2450] = 64'hbd1a7b3d92df5054;
    assign coff[2451] = 64'h8388359be223599e;
    assign coff[2452] = 64'h7c77ca65e223599e;
    assign coff[2453] = 64'h42e584c392df5054;
    assign coff[2454] = 64'he223599e8388359b;
    assign coff[2455] = 64'h92df5054bd1a7b3d;
    assign coff[2456] = 64'h7e6bc8ebebf4fda8;
    assign coff[2457] = 64'h4b387af9986f2d4a;
    assign coff[2458] = 64'hebf4fda881943715;
    assign coff[2459] = 64'h986f2d4ab4c78507;
    assign coff[2460] = 64'h6790d2b6b4c78507;
    assign coff[2461] = 64'h140b025881943715;
    assign coff[2462] = 64'hb4c78507986f2d4a;
    assign coff[2463] = 64'h81943715ebf4fda8;
    assign coff[2464] = 64'h660b91afb2baabde;
    assign coff[2465] = 64'h1184a427813455e6;
    assign coff[2466] = 64'hb2baabde99f46e51;
    assign coff[2467] = 64'h813455e6ee7b5bd9;
    assign coff[2468] = 64'h7ecbaa1aee7b5bd9;
    assign coff[2469] = 64'h4d45542299f46e51;
    assign coff[2470] = 64'hee7b5bd9813455e6;
    assign coff[2471] = 64'h99f46e51b2baabde;
    assign coff[2472] = 64'h7bd9047cdfa97e0f;
    assign coff[2473] = 64'h40b50b46918f60d6;
    assign coff[2474] = 64'hdfa97e0f8426fb84;
    assign coff[2475] = 64'h918f60d6bf4af4ba;
    assign coff[2476] = 64'h6e709f2abf4af4ba;
    assign coff[2477] = 64'h205681f18426fb84;
    assign coff[2478] = 64'hbf4af4ba918f60d6;
    assign coff[2479] = 64'h8426fb84dfa97e0f;
    assign coff[2480] = 64'h7328c1ffc81f3834;
    assign coff[2481] = 64'h29eb0957870ef2f1;
    assign coff[2482] = 64'hc81f38348cd73e01;
    assign coff[2483] = 64'h870ef2f1d614f6a9;
    assign coff[2484] = 64'h78f10d0fd614f6a9;
    assign coff[2485] = 64'h37e0c7cc8cd73e01;
    assign coff[2486] = 64'hd614f6a9870ef2f1;
    assign coff[2487] = 64'h8cd73e01c81f3834;
    assign coff[2488] = 64'h7fc6df08f871e759;
    assign coff[2489] = 64'h5502775ca04e4efc;
    assign coff[2490] = 64'hf871e759803920f8;
    assign coff[2491] = 64'ha04e4efcaafd88a4;
    assign coff[2492] = 64'h5fb1b104aafd88a4;
    assign coff[2493] = 64'h078e18a7803920f8;
    assign coff[2494] = 64'haafd88a4a04e4efc;
    assign coff[2495] = 64'h803920f8f871e759;
    assign coff[2496] = 64'h62217a72add0ad12;
    assign coff[2497] = 64'h0b4684df807f623b;
    assign coff[2498] = 64'hadd0ad129dde858e;
    assign coff[2499] = 64'h807f623bf4b97b21;
    assign coff[2500] = 64'h7f809dc5f4b97b21;
    assign coff[2501] = 64'h522f52ee9dde858e;
    assign coff[2502] = 64'hf4b97b21807f623b;
    assign coff[2503] = 64'h9dde858eadd0ad12;
    assign coff[2504] = 64'h7a1c9eced99fc5d4;
    assign coff[2505] = 64'h3b35d1a58e84a02d;
    assign coff[2506] = 64'hd99fc5d485e36132;
    assign coff[2507] = 64'h8e84a02dc4ca2e5b;
    assign coff[2508] = 64'h717b5fd3c4ca2e5b;
    assign coff[2509] = 64'h26603a2c85e36132;
    assign coff[2510] = 64'hc4ca2e5b8e84a02d;
    assign coff[2511] = 64'h85e36132d99fc5d4;
    assign coff[2512] = 64'h70475839c289e5e7;
    assign coff[2513] = 64'h23eeec788525b228;
    assign coff[2514] = 64'hc289e5e78fb8a7c7;
    assign coff[2515] = 64'h8525b228dc111388;
    assign coff[2516] = 64'h7ada4dd8dc111388;
    assign coff[2517] = 64'h3d761a198fb8a7c7;
    assign coff[2518] = 64'hdc1113888525b228;
    assign coff[2519] = 64'h8fb8a7c7c289e5e7;
    assign coff[2520] = 64'h7f409164f22f2fe1;
    assign coff[2521] = 64'h503635299c3ffbc5;
    assign coff[2522] = 64'hf22f2fe180bf6e9c;
    assign coff[2523] = 64'h9c3ffbc5afc9cad7;
    assign coff[2524] = 64'h63c0043bafc9cad7;
    assign coff[2525] = 64'h0dd0d01f80bf6e9c;
    assign coff[2526] = 64'hafc9cad79c3ffbc5;
    assign coff[2527] = 64'h80bf6e9cf22f2fe1;
    assign coff[2528] = 64'h69b6b9d3b7d45255;
    assign coff[2529] = 64'h17b7f5a382377c4c;
    assign coff[2530] = 64'hb7d452559649462d;
    assign coff[2531] = 64'h82377c4ce8480a5d;
    assign coff[2532] = 64'h7dc883b4e8480a5d;
    assign coff[2533] = 64'h482badab9649462d;
    assign coff[2534] = 64'he8480a5d82377c4c;
    assign coff[2535] = 64'h9649462db7d45255;
    assign coff[2536] = 64'h7d4908d9e5c727dd;
    assign coff[2537] = 64'h460c5cce94de3df8;
    assign coff[2538] = 64'he5c727dd82b6f727;
    assign coff[2539] = 64'h94de3df8b9f3a332;
    assign coff[2540] = 64'h6b21c208b9f3a332;
    assign coff[2541] = 64'h1a38d82382b6f727;
    assign coff[2542] = 64'hb9f3a33294de3df8;
    assign coff[2543] = 64'h82b6f727e5c727dd;
    assign coff[2544] = 64'h75c32634cdd700a4;
    assign coff[2545] = 64'h2fcd4c198942ca39;
    assign coff[2546] = 64'hcdd700a48a3cd9cc;
    assign coff[2547] = 64'h8942ca39d032b3e7;
    assign coff[2548] = 64'h76bd35c7d032b3e7;
    assign coff[2549] = 64'h3228ff5c8a3cd9cc;
    assign coff[2550] = 64'hd032b3e78942ca39;
    assign coff[2551] = 64'h8a3cd9cccdd700a4;
    assign coff[2552] = 64'h7ffe5f03feb947a0;
    assign coff[2553] = 64'h599a4c12a497a693;
    assign coff[2554] = 64'hfeb947a08001a0fd;
    assign coff[2555] = 64'ha497a693a665b3ee;
    assign coff[2556] = 64'h5b68596da665b3ee;
    assign coff[2557] = 64'h0146b8608001a0fd;
    assign coff[2558] = 64'ha665b3eea497a693;
    assign coff[2559] = 64'h8001a0fdfeb947a0;
    assign coff[2560] = 64'h5b452288a641d58c;
    assign coff[2561] = 64'h011474f680012a8e;
    assign coff[2562] = 64'ha641d58ca4badd78;
    assign coff[2563] = 64'h80012a8efeeb8b0a;
    assign coff[2564] = 64'h7ffed572feeb8b0a;
    assign coff[2565] = 64'h59be2a74a4badd78;
    assign coff[2566] = 64'hfeeb8b0a80012a8e;
    assign coff[2567] = 64'ha4badd78a641d58c;
    assign coff[2568] = 64'h76aa670dd00416a3;
    assign coff[2569] = 64'h31fabcbd8a29303b;
    assign coff[2570] = 64'hd00416a3895598f3;
    assign coff[2571] = 64'h8a29303bce054343;
    assign coff[2572] = 64'h75d6cfc5ce054343;
    assign coff[2573] = 64'h2ffbe95d895598f3;
    assign coff[2574] = 64'hce0543438a29303b;
    assign coff[2575] = 64'h895598f3d00416a3;
    assign coff[2576] = 64'h6b0637c1b9c99688;
    assign coff[2577] = 64'h1a07a31182acb4b0;
    assign coff[2578] = 64'hb9c9968894f9c83f;
    assign coff[2579] = 64'h82acb4b0e5f85cef;
    assign coff[2580] = 64'h7d534b50e5f85cef;
    assign coff[2581] = 64'h4636697894f9c83f;
    assign coff[2582] = 64'he5f85cef82acb4b0;
    assign coff[2583] = 64'h94f9c83fb9c99688;
    assign coff[2584] = 64'h7dbf298de816a716;
    assign coff[2585] = 64'h48022499962cf6f2;
    assign coff[2586] = 64'he816a7168240d673;
    assign coff[2587] = 64'h962cf6f2b7fddb67;
    assign coff[2588] = 64'h69d3090eb7fddb67;
    assign coff[2589] = 64'h17e958ea8240d673;
    assign coff[2590] = 64'hb7fddb67962cf6f2;
    assign coff[2591] = 64'h8240d673e816a716;
    assign coff[2592] = 64'h63a07cc7afa2a50f;
    assign coff[2593] = 64'h0d9ed64680ba0b85;
    assign coff[2594] = 64'hafa2a50f9c5f8339;
    assign coff[2595] = 64'h80ba0b85f26129ba;
    assign coff[2596] = 64'h7f45f47bf26129ba;
    assign coff[2597] = 64'h505d5af19c5f8339;
    assign coff[2598] = 64'hf26129ba80ba0b85;
    assign coff[2599] = 64'h9c5f8339afa2a50f;
    assign coff[2600] = 64'h7acc27f7dbe0d7cd;
    assign coff[2601] = 64'h3d49fde18fa08dab;
    assign coff[2602] = 64'hdbe0d7cd8533d809;
    assign coff[2603] = 64'h8fa08dabc2b6021f;
    assign coff[2604] = 64'h705f7255c2b6021f;
    assign coff[2605] = 64'h241f28338533d809;
    assign coff[2606] = 64'hc2b6021f8fa08dab;
    assign coff[2607] = 64'h8533d809dbe0d7cd;
    assign coff[2608] = 64'h7164169dc49da27a;
    assign coff[2609] = 64'h2630433385d458a6;
    assign coff[2610] = 64'hc49da27a8e9be963;
    assign coff[2611] = 64'h85d458a6d9cfbccd;
    assign coff[2612] = 64'h7a2ba75ad9cfbccd;
    assign coff[2613] = 64'h3b625d868e9be963;
    assign coff[2614] = 64'hd9cfbccd85d458a6;
    assign coff[2615] = 64'h8e9be963c49da27a;
    assign coff[2616] = 64'h7f7c2668f4876a10;
    assign coff[2617] = 64'h5208c36a9dbe4701;
    assign coff[2618] = 64'hf4876a108083d998;
    assign coff[2619] = 64'h9dbe4701adf73c96;
    assign coff[2620] = 64'h6241b8ffadf73c96;
    assign coff[2621] = 64'h0b7895f08083d998;
    assign coff[2622] = 64'hadf73c969dbe4701;
    assign coff[2623] = 64'h8083d998f4876a10;
    assign coff[2624] = 64'h5f90478aaad7fafb;
    assign coff[2625] = 64'h075bea8c8036334e;
    assign coff[2626] = 64'haad7fafba06fb876;
    assign coff[2627] = 64'h8036334ef8a41574;
    assign coff[2628] = 64'h7fc9ccb2f8a41574;
    assign coff[2629] = 64'h55280505a06fb876;
    assign coff[2630] = 64'hf8a415748036334e;
    assign coff[2631] = 64'ha06fb876aad7fafb;
    assign coff[2632] = 64'h78e08dabd5e57b85;
    assign coff[2633] = 64'h37b38a6d8cc1556a;
    assign coff[2634] = 64'hd5e57b85871f7255;
    assign coff[2635] = 64'h8cc1556ac84c7593;
    assign coff[2636] = 64'h733eaa96c84c7593;
    assign coff[2637] = 64'h2a1a847b871f7255;
    assign coff[2638] = 64'hc84c75938cc1556a;
    assign coff[2639] = 64'h871f7255d5e57b85;
    assign coff[2640] = 64'h6e572d93bf1f9b16;
    assign coff[2641] = 64'h2025dcec841a521a;
    assign coff[2642] = 64'hbf1f9b1691a8d26d;
    assign coff[2643] = 64'h841a521adfda2314;
    assign coff[2644] = 64'h7be5ade6dfda2314;
    assign coff[2645] = 64'h40e064ea91a8d26d;
    assign coff[2646] = 64'hdfda2314841a521a;
    assign coff[2647] = 64'h91a8d26dbf1f9b16;
    assign coff[2648] = 64'h7ec4bf36ee499253;
    assign coff[2649] = 64'h4d1d3b7a99d61e14;
    assign coff[2650] = 64'hee499253813b40ca;
    assign coff[2651] = 64'h99d61e14b2e2c486;
    assign coff[2652] = 64'h6629e1ecb2e2c486;
    assign coff[2653] = 64'h11b66dad813b40ca;
    assign coff[2654] = 64'hb2e2c48699d61e14;
    assign coff[2655] = 64'h813b40caee499253;
    assign coff[2656] = 64'h677340bab49edf45;
    assign coff[2657] = 64'h13d95b93818c61e3;
    assign coff[2658] = 64'hb49edf45988cbf46;
    assign coff[2659] = 64'h818c61e3ec26a46d;
    assign coff[2660] = 64'h7e739e1dec26a46d;
    assign coff[2661] = 64'h4b6120bb988cbf46;
    assign coff[2662] = 64'hec26a46d818c61e3;
    assign coff[2663] = 64'h988cbf46b49edf45;
    assign coff[2664] = 64'h7c6c06c0e1f27b0b;
    assign coff[2665] = 64'h42baa4e692c51392;
    assign coff[2666] = 64'he1f27b0b8393f940;
    assign coff[2667] = 64'h92c51392bd455b1a;
    assign coff[2668] = 64'h6d3aec6ebd455b1a;
    assign coff[2669] = 64'h1e0d84f58393f940;
    assign coff[2670] = 64'hbd455b1a92c51392;
    assign coff[2671] = 64'h8393f940e1f27b0b;
    assign coff[2672] = 64'h742b1144ca404992;
    assign coff[2673] = 64'h2c231c3387d9b7b7;
    assign coff[2674] = 64'hca4049928bd4eebc;
    assign coff[2675] = 64'h87d9b7b7d3dce3cd;
    assign coff[2676] = 64'h78264849d3dce3cd;
    assign coff[2677] = 64'h35bfb66e8bd4eebc;
    assign coff[2678] = 64'hd3dce3cd87d9b7b7;
    assign coff[2679] = 64'h8bd4eebcca404992;
    assign coff[2680] = 64'h7fe4ee06facc54e0;
    assign coff[2681] = 64'h56c1b3a1a1e308e4;
    assign coff[2682] = 64'hfacc54e0801b11fa;
    assign coff[2683] = 64'ha1e308e4a93e4c5f;
    assign coff[2684] = 64'h5e1cf71ca93e4c5f;
    assign coff[2685] = 64'h0533ab20801b11fa;
    assign coff[2686] = 64'ha93e4c5fa1e308e4;
    assign coff[2687] = 64'h801b11fafacc54e0;
    assign coff[2688] = 64'h5d71e979a88629a5;
    assign coff[2689] = 64'h043883108011d1d0;
    assign coff[2690] = 64'ha88629a5a28e1687;
    assign coff[2691] = 64'h8011d1d0fbc77cf0;
    assign coff[2692] = 64'h7fee2e30fbc77cf0;
    assign coff[2693] = 64'h5779d65ba28e1687;
    assign coff[2694] = 64'hfbc77cf08011d1d0;
    assign coff[2695] = 64'ha28e1687a88629a5;
    assign coff[2696] = 64'h77ceb725d2f14fba;
    assign coff[2697] = 64'h34db36df8b6c45cc;
    assign coff[2698] = 64'hd2f14fba883148db;
    assign coff[2699] = 64'h8b6c45cccb24c921;
    assign coff[2700] = 64'h7493ba34cb24c921;
    assign coff[2701] = 64'h2d0eb046883148db;
    assign coff[2702] = 64'hcb24c9218b6c45cc;
    assign coff[2703] = 64'h883148dbd2f14fba;
    assign coff[2704] = 64'h6cb71482bc6f6333;
    assign coff[2705] = 64'h1d18fe548359e70d;
    assign coff[2706] = 64'hbc6f63339348eb7e;
    assign coff[2707] = 64'h8359e70de2e701ac;
    assign coff[2708] = 64'h7ca618f3e2e701ac;
    assign coff[2709] = 64'h43909ccd9348eb7e;
    assign coff[2710] = 64'he2e701ac8359e70d;
    assign coff[2711] = 64'h9348eb7ebc6f6333;
    assign coff[2712] = 64'h7e4bb13ceb2e81ca;
    assign coff[2713] = 64'h4a95703097f9853d;
    assign coff[2714] = 64'heb2e81ca81b44ec4;
    assign coff[2715] = 64'h97f9853db56a8fd0;
    assign coff[2716] = 64'h68067ac3b56a8fd0;
    assign coff[2717] = 64'h14d17e3681b44ec4;
    assign coff[2718] = 64'hb56a8fd097f9853d;
    assign coff[2719] = 64'h81b44ec4eb2e81ca;
    assign coff[2720] = 64'h6591b38cb21ac0a6;
    assign coff[2721] = 64'h10bd635681196de9;
    assign coff[2722] = 64'hb21ac0a69a6e4c74;
    assign coff[2723] = 64'h81196de9ef429caa;
    assign coff[2724] = 64'h7ee69217ef429caa;
    assign coff[2725] = 64'h4de53f5a9a6e4c74;
    assign coff[2726] = 64'hef429caa81196de9;
    assign coff[2727] = 64'h9a6e4c74b21ac0a6;
    assign coff[2728] = 64'h7ba59feedee71c24;
    assign coff[2729] = 64'h40074132912a44f0;
    assign coff[2730] = 64'hdee71c24845a6012;
    assign coff[2731] = 64'h912a44f0bff8bece;
    assign coff[2732] = 64'h6ed5bb10bff8bece;
    assign coff[2733] = 64'h2118e3dc845a6012;
    assign coff[2734] = 64'hbff8bece912a44f0;
    assign coff[2735] = 64'h845a6012dee71c24;
    assign coff[2736] = 64'h72d06e2bc76a992a;
    assign coff[2737] = 64'h292cdc6d86cdaffa;
    assign coff[2738] = 64'hc76a992a8d2f91d5;
    assign coff[2739] = 64'h86cdaffad6d32393;
    assign coff[2740] = 64'h79325006d6d32393;
    assign coff[2741] = 64'h389566d68d2f91d5;
    assign coff[2742] = 64'hd6d3239386cdaffa;
    assign coff[2743] = 64'h8d2f91d5c76a992a;
    assign coff[2744] = 64'h7fba6357f7a93ae0;
    assign coff[2745] = 64'h546bbdd79fc93cdb;
    assign coff[2746] = 64'hf7a93ae080459ca9;
    assign coff[2747] = 64'h9fc93cdbab944229;
    assign coff[2748] = 64'h6036c325ab944229;
    assign coff[2749] = 64'h0856c52080459ca9;
    assign coff[2750] = 64'hab9442299fc93cdb;
    assign coff[2751] = 64'h80459ca9f7a93ae0;
    assign coff[2752] = 64'h619fe918ad36edfc;
    assign coff[2753] = 64'h0a7e2f85806e496c;
    assign coff[2754] = 64'had36edfc9e6016e8;
    assign coff[2755] = 64'h806e496cf581d07b;
    assign coff[2756] = 64'h7f91b694f581d07b;
    assign coff[2757] = 64'h52c912049e6016e8;
    assign coff[2758] = 64'hf581d07b806e496c;
    assign coff[2759] = 64'h9e6016e8ad36edfc;
    assign coff[2760] = 64'h79dfc064d8e0256a;
    assign coff[2761] = 64'h3a8347178e282a7b;
    assign coff[2762] = 64'hd8e0256a86203f9c;
    assign coff[2763] = 64'h8e282a7bc57cb8e9;
    assign coff[2764] = 64'h71d7d585c57cb8e9;
    assign coff[2765] = 64'h271fda9686203f9c;
    assign coff[2766] = 64'hc57cb8e98e282a7b;
    assign coff[2767] = 64'h86203f9cd8e0256a;
    assign coff[2768] = 64'h6fe642cac1d9d412;
    assign coff[2769] = 64'h232dc66d84edd82d;
    assign coff[2770] = 64'hc1d9d4129019bd36;
    assign coff[2771] = 64'h84edd82ddcd23993;
    assign coff[2772] = 64'h7b1227d3dcd23993;
    assign coff[2773] = 64'h3e262bee9019bd36;
    assign coff[2774] = 64'hdcd2399384edd82d;
    assign coff[2775] = 64'h9019bd36c1d9d412;
    assign coff[2776] = 64'h7f2a40d2f1675e17;
    assign coff[2777] = 64'h4f9922939bc277fa;
    assign coff[2778] = 64'hf1675e1780d5bf2e;
    assign coff[2779] = 64'h9bc277fab066dd6d;
    assign coff[2780] = 64'h643d8806b066dd6d;
    assign coff[2781] = 64'h0e98a1e980d5bf2e;
    assign coff[2782] = 64'hb066dd6d9bc277fa;
    assign coff[2783] = 64'h80d5bf2ef1675e17;
    assign coff[2784] = 64'h6944da10b72e9d9b;
    assign coff[2785] = 64'h16f2443e8212d5b9;
    assign coff[2786] = 64'hb72e9d9b96bb25f0;
    assign coff[2787] = 64'h8212d5b9e90dbbc2;
    assign coff[2788] = 64'h7ded2a47e90dbbc2;
    assign coff[2789] = 64'h48d1626596bb25f0;
    assign coff[2790] = 64'he90dbbc28212d5b9;
    assign coff[2791] = 64'h96bb25f0b72e9d9b;
    assign coff[2792] = 64'h7d1f3dd6e5027c53;
    assign coff[2793] = 64'h4563be609470ba39;
    assign coff[2794] = 64'he5027c5382e0c22a;
    assign coff[2795] = 64'h9470ba39ba9c41a0;
    assign coff[2796] = 64'h6b8f45c7ba9c41a0;
    assign coff[2797] = 64'h1afd83ad82e0c22a;
    assign coff[2798] = 64'hba9c41a09470ba39;
    assign coff[2799] = 64'h82e0c22ae5027c53;
    assign coff[2800] = 64'h7573ca75cd1e43ca;
    assign coff[2801] = 64'h2f128d9988f84687;
    assign coff[2802] = 64'hcd1e43ca8a8c358b;
    assign coff[2803] = 64'h88f84687d0ed7267;
    assign coff[2804] = 64'h7707b979d0ed7267;
    assign coff[2805] = 64'h32e1bc368a8c358b;
    assign coff[2806] = 64'hd0ed726788f84687;
    assign coff[2807] = 64'h8a8c358bcd1e43ca;
    assign coff[2808] = 64'h7ffbbfe6fdf03c3a;
    assign coff[2809] = 64'h590a4893a40b582e;
    assign coff[2810] = 64'hfdf03c3a8004401a;
    assign coff[2811] = 64'ha40b582ea6f5b76d;
    assign coff[2812] = 64'h5bf4a7d2a6f5b76d;
    assign coff[2813] = 64'h020fc3c68004401a;
    assign coff[2814] = 64'ha6f5b76da40b582e;
    assign coff[2815] = 64'h8004401afdf03c3a;
    assign coff[2816] = 64'h5c5d4dcca7624a4d;
    assign coff[2817] = 64'h02a68917800706ac;
    assign coff[2818] = 64'ha7624a4da3a2b234;
    assign coff[2819] = 64'h800706acfd5976e9;
    assign coff[2820] = 64'h7ff8f954fd5976e9;
    assign coff[2821] = 64'h589db5b3a3a2b234;
    assign coff[2822] = 64'hfd5976e9800706ac;
    assign coff[2823] = 64'ha3a2b234a7624a4d;
    assign coff[2824] = 64'h773edb8bd179cd99;
    assign coff[2825] = 64'h336bf78f8ac87894;
    assign coff[2826] = 64'hd179cd9988c12475;
    assign coff[2827] = 64'h8ac87894cc940871;
    assign coff[2828] = 64'h7537876ccc940871;
    assign coff[2829] = 64'h2e86326788c12475;
    assign coff[2830] = 64'hcc9408718ac87894;
    assign coff[2831] = 64'h88c12475d179cd99;
    assign coff[2832] = 64'h6be0ba7bbb1b28e4;
    assign coff[2833] = 64'h1b90d8bb8300e50b;
    assign coff[2834] = 64'hbb1b28e4941f4585;
    assign coff[2835] = 64'h8300e50be46f2745;
    assign coff[2836] = 64'h7cff1af5e46f2745;
    assign coff[2837] = 64'h44e4d71c941f4585;
    assign coff[2838] = 64'he46f27458300e50b;
    assign coff[2839] = 64'h941f4585bb1b28e4;
    assign coff[2840] = 64'h7e07db52e9a22610;
    assign coff[2841] = 64'h494d341e97113847;
    assign coff[2842] = 64'he9a2261081f824ae;
    assign coff[2843] = 64'h97113847b6b2cbe2;
    assign coff[2844] = 64'h68eec7b9b6b2cbe2;
    assign coff[2845] = 64'h165dd9f081f824ae;
    assign coff[2846] = 64'hb6b2cbe297113847;
    assign coff[2847] = 64'h81f824aee9a22610;
    assign coff[2848] = 64'h649b08a0b0dd2c56;
    assign coff[2849] = 64'h0f2e67b880e74987;
    assign coff[2850] = 64'hb0dd2c569b64f760;
    assign coff[2851] = 64'h80e74987f0d19848;
    assign coff[2852] = 64'h7f18b679f0d19848;
    assign coff[2853] = 64'h4f22d3aa9b64f760;
    assign coff[2854] = 64'hf0d1984880e74987;
    assign coff[2855] = 64'h9b64f760b0dd2c56;
    assign coff[2856] = 64'h7b3b4410dd634f2b;
    assign coff[2857] = 64'h3ea9d4c390634287;
    assign coff[2858] = 64'hdd634f2b84c4bbf0;
    assign coff[2859] = 64'h90634287c1562b3d;
    assign coff[2860] = 64'h6f9cbd79c1562b3d;
    assign coff[2861] = 64'h229cb0d584c4bbf0;
    assign coff[2862] = 64'hc1562b3d90634287;
    assign coff[2863] = 64'h84c4bbf0dd634f2b;
    assign coff[2864] = 64'h721c7580c602ffaa;
    assign coff[2865] = 64'h27af53a6864eabcb;
    assign coff[2866] = 64'hc602ffaa8de38a80;
    assign coff[2867] = 64'h864eabcbd850ac5a;
    assign coff[2868] = 64'h79b15435d850ac5a;
    assign coff[2869] = 64'h39fd00568de38a80;
    assign coff[2870] = 64'hd850ac5a864eabcb;
    assign coff[2871] = 64'h8de38a80c602ffaa;
    assign coff[2872] = 64'h7f9dbaa0f6182196;
    assign coff[2873] = 64'h533bdb5d9ec1e210;
    assign coff[2874] = 64'hf618219680624560;
    assign coff[2875] = 64'h9ec1e210acc424a3;
    assign coff[2876] = 64'h613e1df0acc424a3;
    assign coff[2877] = 64'h09e7de6a80624560;
    assign coff[2878] = 64'hacc424a39ec1e210;
    assign coff[2879] = 64'h80624560f6182196;
    assign coff[2880] = 64'h6099f505ac05d613;
    assign coff[2881] = 64'h08ed3916804fc841;
    assign coff[2882] = 64'hac05d6139f660afb;
    assign coff[2883] = 64'h804fc841f712c6ea;
    assign coff[2884] = 64'h7fb037bff712c6ea;
    assign coff[2885] = 64'h53fa29ed9f660afb;
    assign coff[2886] = 64'hf712c6ea804fc841;
    assign coff[2887] = 64'h9f660afbac05d613;
    assign coff[2888] = 64'h79627e08d7620808;
    assign coff[2889] = 64'h391c82978d728aa9;
    assign coff[2890] = 64'hd7620808869d81f8;
    assign coff[2891] = 64'h8d728aa9c6e37d69;
    assign coff[2892] = 64'h728d7557c6e37d69;
    assign coff[2893] = 64'h289df7f8869d81f8;
    assign coff[2894] = 64'hc6e37d698d728aa9;
    assign coff[2895] = 64'h869d81f8d7620808;
    assign coff[2896] = 64'h6f20dc92c07b7e23;
    assign coff[2897] = 64'h21aa77cf8481b3bb;
    assign coff[2898] = 64'hc07b7e2390df236e;
    assign coff[2899] = 64'h8481b3bbde558831;
    assign coff[2900] = 64'h7b7e4c45de558831;
    assign coff[2901] = 64'h3f8481dd90df236e;
    assign coff[2902] = 64'hde5588318481b3bb;
    assign coff[2903] = 64'h90df236ec07b7e23;
    assign coff[2904] = 64'h7ef9f29defd8287c;
    assign coff[2905] = 64'h4e5cb1b99aca5795;
    assign coff[2906] = 64'hefd8287c81060d63;
    assign coff[2907] = 64'h9aca5795b1a34e47;
    assign coff[2908] = 64'h6535a86bb1a34e47;
    assign coff[2909] = 64'h1027d78481060d63;
    assign coff[2910] = 64'hb1a34e479aca5795;
    assign coff[2911] = 64'h81060d63efd8287c;
    assign coff[2912] = 64'h685e106cb5e550c1;
    assign coff[2913] = 64'h1566398281cd2d0c;
    assign coff[2914] = 64'hb5e550c197a1ef94;
    assign coff[2915] = 64'h81cd2d0cea99c67e;
    assign coff[2916] = 64'h7e32d2f4ea99c67e;
    assign coff[2917] = 64'h4a1aaf3f97a1ef94;
    assign coff[2918] = 64'hea99c67e81cd2d0c;
    assign coff[2919] = 64'h97a1ef94b5e550c1;
    assign coff[2920] = 64'h7cc80a0fe379eeed;
    assign coff[2921] = 64'h441081849398cff5;
    assign coff[2922] = 64'he379eeed8337f5f1;
    assign coff[2923] = 64'h9398cff5bbef7e7c;
    assign coff[2924] = 64'h6c67300bbbef7e7c;
    assign coff[2925] = 64'h1c8611138337f5f1;
    assign coff[2926] = 64'hbbef7e7c9398cff5;
    assign coff[2927] = 64'h8337f5f1e379eeed;
    assign coff[2928] = 64'h74d1ae55cbae447f;
    assign coff[2929] = 64'h2d9bb5f68866b0ef;
    assign coff[2930] = 64'hcbae447f8b2e51ab;
    assign coff[2931] = 64'h8866b0efd2644a0a;
    assign coff[2932] = 64'h77994f11d2644a0a;
    assign coff[2933] = 64'h3451bb818b2e51ab;
    assign coff[2934] = 64'hd2644a0a8866b0ef;
    assign coff[2935] = 64'h8b2e51abcbae447f;
    assign coff[2936] = 64'h7ff2ce5bfc5e36a0;
    assign coff[2937] = 64'h57e7afe4a2f56566;
    assign coff[2938] = 64'hfc5e36a0800d31a5;
    assign coff[2939] = 64'ha2f56566a818501c;
    assign coff[2940] = 64'h5d0a9a9aa818501c;
    assign coff[2941] = 64'h03a1c960800d31a5;
    assign coff[2942] = 64'ha818501ca2f56566;
    assign coff[2943] = 64'h800d31a5fc5e36a0;
    assign coff[2944] = 64'h5e82eae5a9ad6855;
    assign coff[2945] = 64'h05ca536180218b8f;
    assign coff[2946] = 64'ha9ad6855a17d151b;
    assign coff[2947] = 64'h80218b8ffa35ac9f;
    assign coff[2948] = 64'h7fde7471fa35ac9f;
    assign coff[2949] = 64'h565297aba17d151b;
    assign coff[2950] = 64'hfa35ac9f80218b8f;
    assign coff[2951] = 64'ha17d151ba9ad6855;
    assign coff[2952] = 64'h7859f44fd46a8e8d;
    assign coff[2953] = 64'h36486c868c149192;
    assign coff[2954] = 64'hd46a8e8d87a60bb1;
    assign coff[2955] = 64'h8c149192c9b7937a;
    assign coff[2956] = 64'h73eb6e6ec9b7937a;
    assign coff[2957] = 64'h2b95717387a60bb1;
    assign coff[2958] = 64'hc9b7937a8c149192;
    assign coff[2959] = 64'h87a60bb1d46a8e8d;
    assign coff[2960] = 64'h6d893d93bdc63856;
    assign coff[2961] = 64'h1ea004c183b7b746;
    assign coff[2962] = 64'hbdc638569276c26d;
    assign coff[2963] = 64'h83b7b746e15ffb3f;
    assign coff[2964] = 64'h7c4848bae15ffb3f;
    assign coff[2965] = 64'h4239c7aa9276c26d;
    assign coff[2966] = 64'he15ffb3f83b7b746;
    assign coff[2967] = 64'h9276c26dbdc63856;
    assign coff[2968] = 64'h7e8aa8acecbbaafb;
    assign coff[2969] = 64'h4bdacc2898e5d4e0;
    assign coff[2970] = 64'hecbbaafb81755754;
    assign coff[2971] = 64'h98e5d4e0b42533d8;
    assign coff[2972] = 64'h671a2b20b42533d8;
    assign coff[2973] = 64'h1344550581755754;
    assign coff[2974] = 64'hb42533d898e5d4e0;
    assign coff[2975] = 64'h81755754ecbbaafb;
    assign coff[2976] = 64'h66847408b35b55bf;
    assign coff[2977] = 64'h124bb9be815076bd;
    assign coff[2978] = 64'hb35b55bf997b8bf8;
    assign coff[2979] = 64'h815076bdedb44642;
    assign coff[2980] = 64'h7eaf8943edb44642;
    assign coff[2981] = 64'h4ca4aa41997b8bf8;
    assign coff[2982] = 64'hedb44642815076bd;
    assign coff[2983] = 64'h997b8bf8b35b55bf;
    assign coff[2984] = 64'h7c0b3777e06c2fc4;
    assign coff[2985] = 64'h416235b291f58d3b;
    assign coff[2986] = 64'he06c2fc483f4c889;
    assign coff[2987] = 64'h91f58d3bbe9dca4e;
    assign coff[2988] = 64'h6e0a72c5be9dca4e;
    assign coff[2989] = 64'h1f93d03c83f4c889;
    assign coff[2990] = 64'hbe9dca4e91f58d3b;
    assign coff[2991] = 64'h83f4c889e06c2fc4;
    assign coff[2992] = 64'h737ff9aec8d4611d;
    assign coff[2993] = 64'h2aa8ced387516050;
    assign coff[2994] = 64'hc8d4611d8c800652;
    assign coff[2995] = 64'h87516050d557312d;
    assign coff[2996] = 64'h78ae9fb0d557312d;
    assign coff[2997] = 64'h372b9ee38c800652;
    assign coff[2998] = 64'hd557312d87516050;
    assign coff[2999] = 64'h8c800652c8d4611d;
    assign coff[3000] = 64'h7fd21f72f93aa676;
    assign coff[3001] = 64'h55985f20a0d44d3b;
    assign coff[3002] = 64'hf93aa676802de08e;
    assign coff[3003] = 64'ha0d44d3baa67a0e0;
    assign coff[3004] = 64'h5f2bb2c5aa67a0e0;
    assign coff[3005] = 64'h06c5598a802de08e;
    assign coff[3006] = 64'haa67a0e0a0d44d3b;
    assign coff[3007] = 64'h802de08ef93aa676;
    assign coff[3008] = 64'h62a219aaae6b36f0;
    assign coff[3009] = 64'h0c0ebe668091b5a2;
    assign coff[3010] = 64'hae6b36f09d5de656;
    assign coff[3011] = 64'h8091b5a2f3f1419a;
    assign coff[3012] = 64'h7f6e4a5ef3f1419a;
    assign coff[3013] = 64'h5194c9109d5de656;
    assign coff[3014] = 64'hf3f1419a8091b5a2;
    assign coff[3015] = 64'h9d5de656ae6b36f0;
    assign coff[3016] = 64'h7a584febda5fc4ef;
    assign coff[3017] = 64'h3be7ca1a8ee22de0;
    assign coff[3018] = 64'hda5fc4ef85a7b015;
    assign coff[3019] = 64'h8ee22de0c41835e6;
    assign coff[3020] = 64'h711dd220c41835e6;
    assign coff[3021] = 64'h25a03b1185a7b015;
    assign coff[3022] = 64'hc41835e68ee22de0;
    assign coff[3023] = 64'h85a7b015da5fc4ef;
    assign coff[3024] = 64'h70a7589fc33a8f62;
    assign coff[3025] = 64'h24afb9da855ebb44;
    assign coff[3026] = 64'hc33a8f628f58a761;
    assign coff[3027] = 64'h855ebb44db504626;
    assign coff[3028] = 64'h7aa144bcdb504626;
    assign coff[3029] = 64'h3cc5709e8f58a761;
    assign coff[3030] = 64'hdb504626855ebb44;
    assign coff[3031] = 64'h8f58a761c33a8f62;
    assign coff[3032] = 64'h7f55a7faf2f723c1;
    assign coff[3033] = 64'h50d281d59cbe75b0;
    assign coff[3034] = 64'hf2f723c180aa5806;
    assign coff[3035] = 64'h9cbe75b0af2d7e2b;
    assign coff[3036] = 64'h63418a50af2d7e2b;
    assign coff[3037] = 64'h0d08dc3f80aa5806;
    assign coff[3038] = 64'haf2d7e2b9cbe75b0;
    assign coff[3039] = 64'h80aa5806f2f723c1;
    assign coff[3040] = 64'h6a2794c1b87ab922;
    assign coff[3041] = 64'h187d6c82825d593a;
    assign coff[3042] = 64'hb87ab92295d86b3f;
    assign coff[3043] = 64'h825d593ae782937e;
    assign coff[3044] = 64'h7da2a6c6e782937e;
    assign coff[3045] = 64'h478546de95d86b3f;
    assign coff[3046] = 64'he782937e825d593a;
    assign coff[3047] = 64'h95d86b3fb87ab922;
    assign coff[3048] = 64'h7d719ebae68c141a;
    assign coff[3049] = 64'h46b44e65954cca0c;
    assign coff[3050] = 64'he68c141a828e6146;
    assign coff[3051] = 64'h954cca0cb94bb19b;
    assign coff[3052] = 64'h6ab335f4b94bb19b;
    assign coff[3053] = 64'h1973ebe6828e6146;
    assign coff[3054] = 64'hb94bb19b954cca0c;
    assign coff[3055] = 64'h828e6146e68c141a;
    assign coff[3056] = 64'h76115f63ce903942;
    assign coff[3057] = 64'h308794a6898e72e4;
    assign coff[3058] = 64'hce90394289eea09d;
    assign coff[3059] = 64'h898e72e4cf786b5a;
    assign coff[3060] = 64'h76718d1ccf786b5a;
    assign coff[3061] = 64'h316fc6be89eea09d;
    assign coff[3062] = 64'hcf786b5a898e72e4;
    assign coff[3063] = 64'h89eea09dce903942;
    assign coff[3064] = 64'h7fffc251ff82562c;
    assign coff[3065] = 64'h5a29727ba524d683;
    assign coff[3066] = 64'hff82562c80003daf;
    assign coff[3067] = 64'ha524d683a5d68d85;
    assign coff[3068] = 64'h5adb297da5d68d85;
    assign coff[3069] = 64'h007da9d480003daf;
    assign coff[3070] = 64'ha5d68d85a524d683;
    assign coff[3071] = 64'h80003dafff82562c;
    assign coff[3072] = 64'h5afe8a8ba5fa4252;
    assign coff[3073] = 64'h00afeda8800078e7;
    assign coff[3074] = 64'ha5fa4252a5017575;
    assign coff[3075] = 64'h800078e7ff501258;
    assign coff[3076] = 64'h7fff8719ff501258;
    assign coff[3077] = 64'h5a05bdaea5017575;
    assign coff[3078] = 64'hff501258800078e7;
    assign coff[3079] = 64'ha5017575a5fa4252;
    assign coff[3080] = 64'h768492b4cfa6f255;
    assign coff[3081] = 64'h319e20678a0213a0;
    assign coff[3082] = 64'hcfa6f255897b6d4c;
    assign coff[3083] = 64'h8a0213a0ce61df99;
    assign coff[3084] = 64'h75fdec60ce61df99;
    assign coff[3085] = 64'h30590dab897b6d4c;
    assign coff[3086] = 64'hce61df998a0213a0;
    assign coff[3087] = 64'h897b6d4ccfa6f255;
    assign coff[3088] = 64'h6acef1b2b9759db6;
    assign coff[3089] = 64'h19a52ceb829869be;
    assign coff[3090] = 64'hb9759db695310e4e;
    assign coff[3091] = 64'h829869bee65ad315;
    assign coff[3092] = 64'h7d679642e65ad315;
    assign coff[3093] = 64'h468a624a95310e4e;
    assign coff[3094] = 64'he65ad315829869be;
    assign coff[3095] = 64'h95310e4eb9759db6;
    assign coff[3096] = 64'h7dac3b15e7b3eb9f;
    assign coff[3097] = 64'h47aef12c95f48977;
    assign coff[3098] = 64'he7b3eb9f8253c4eb;
    assign coff[3099] = 64'h95f48977b8510ed4;
    assign coff[3100] = 64'h6a0b7689b8510ed4;
    assign coff[3101] = 64'h184c14618253c4eb;
    assign coff[3102] = 64'hb8510ed495f48977;
    assign coff[3103] = 64'h8253c4ebe7b3eb9f;
    assign coff[3104] = 64'h63613fcdaf547eb3;
    assign coff[3105] = 64'h0d3adc4e80af8039;
    assign coff[3106] = 64'haf547eb39c9ec033;
    assign coff[3107] = 64'h80af8039f2c523b2;
    assign coff[3108] = 64'h7f507fc7f2c523b2;
    assign coff[3109] = 64'h50ab814d9c9ec033;
    assign coff[3110] = 64'hf2c523b280af8039;
    assign coff[3111] = 64'h9c9ec033af547eb3;
    assign coff[3112] = 64'h7aafa367db807114;
    assign coff[3113] = 64'h3cf1a91c8f708d75;
    assign coff[3114] = 64'hdb80711485505c99;
    assign coff[3115] = 64'h8f708d75c30e56e4;
    assign coff[3116] = 64'h708f728bc30e56e4;
    assign coff[3117] = 64'h247f8eec85505c99;
    assign coff[3118] = 64'hc30e56e48f708d75;
    assign coff[3119] = 64'h85505c99db807114;
    assign coff[3120] = 64'h71354fc0c444a639;
    assign coff[3121] = 64'h25d0439f85b68015;
    assign coff[3122] = 64'hc444a6398ecab040;
    assign coff[3123] = 64'h85b68015da2fbc61;
    assign coff[3124] = 64'h7a497febda2fbc61;
    assign coff[3125] = 64'h3bbb59c78ecab040;
    assign coff[3126] = 64'hda2fbc6185b68015;
    assign coff[3127] = 64'h8ecab040c444a639;
    assign coff[3128] = 64'h7f72fcb4f4234d45;
    assign coff[3129] = 64'h51bb7e759d7df75f;
    assign coff[3130] = 64'hf4234d45808d034c;
    assign coff[3131] = 64'h9d7df75fae44818b;
    assign coff[3132] = 64'h628208a1ae44818b;
    assign coff[3133] = 64'h0bdcb2bb808d034c;
    assign coff[3134] = 64'hae44818b9d7df75f;
    assign coff[3135] = 64'h808d034cf4234d45;
    assign coff[3136] = 64'h5f4d4865aa8d0713;
    assign coff[3137] = 64'h06f78af680309318;
    assign coff[3138] = 64'haa8d0713a0b2b79b;
    assign coff[3139] = 64'h80309318f908750a;
    assign coff[3140] = 64'h7fcf6ce8f908750a;
    assign coff[3141] = 64'h5572f8eda0b2b79b;
    assign coff[3142] = 64'hf908750a80309318;
    assign coff[3143] = 64'ha0b2b79baa8d0713;
    assign coff[3144] = 64'h78bf56f9d58698c0;
    assign coff[3145] = 64'h3758f5f28c95b98f;
    assign coff[3146] = 64'hd58698c08740a907;
    assign coff[3147] = 64'h8c95b98fc8a70a0e;
    assign coff[3148] = 64'h736a4671c8a70a0e;
    assign coff[3149] = 64'h2a7967408740a907;
    assign coff[3150] = 64'hc8a70a0e8c95b98f;
    assign coff[3151] = 64'h8740a907d58698c0;
    assign coff[3152] = 64'h6e24175cbec905d9;
    assign coff[3153] = 64'h1fc4840a8401389b;
    assign coff[3154] = 64'hbec905d991dbe8a4;
    assign coff[3155] = 64'h8401389be03b7bf6;
    assign coff[3156] = 64'h7bfec765e03b7bf6;
    assign coff[3157] = 64'h4136fa2791dbe8a4;
    assign coff[3158] = 64'he03b7bf68401389b;
    assign coff[3159] = 64'h91dbe8a4bec905d9;
    assign coff[3160] = 64'h7eb6aecaede60780;
    assign coff[3161] = 64'h4ccce6849999ace3;
    assign coff[3162] = 64'hede6078081495136;
    assign coff[3163] = 64'h9999ace3b333197c;
    assign coff[3164] = 64'h6666531db333197c;
    assign coff[3165] = 64'h1219f88081495136;
    assign coff[3166] = 64'hb333197c9999ace3;
    assign coff[3167] = 64'h81495136ede60780;
    assign coff[3168] = 64'h6737eceab44db6a8;
    assign coff[3169] = 64'h137604e2817cf201;
    assign coff[3170] = 64'hb44db6a898c81316;
    assign coff[3171] = 64'h817cf201ec89fb1e;
    assign coff[3172] = 64'h7e830dffec89fb1e;
    assign coff[3173] = 64'h4bb2495898c81316;
    assign coff[3174] = 64'hec89fb1e817cf201;
    assign coff[3175] = 64'h98c81316b44db6a8;
    assign coff[3176] = 64'h7c5445e9e190cbd4;
    assign coff[3177] = 64'h4264c6539290cc9b;
    assign coff[3178] = 64'he190cbd483abba17;
    assign coff[3179] = 64'h9290cc9bbd9b39ad;
    assign coff[3180] = 64'h6d6f3365bd9b39ad;
    assign coff[3181] = 64'h1e6f342c83abba17;
    assign coff[3182] = 64'hbd9b39ad9290cc9b;
    assign coff[3183] = 64'h83abba17e190cbd4;
    assign coff[3184] = 64'h7400b69ac9e51d2d;
    assign coff[3185] = 64'h2bc4b12087b7327d;
    assign coff[3186] = 64'hc9e51d2d8bff4966;
    assign coff[3187] = 64'h87b7327dd43b4ee0;
    assign coff[3188] = 64'h7848cd83d43b4ee0;
    assign coff[3189] = 64'h361ae2d38bff4966;
    assign coff[3190] = 64'hd43b4ee087b7327d;
    assign coff[3191] = 64'h8bff4966c9e51d2d;
    assign coff[3192] = 64'h7fe0b0b1fa67e3da;
    assign coff[3193] = 64'h5677ae54a19f027c;
    assign coff[3194] = 64'hfa67e3da801f4f4f;
    assign coff[3195] = 64'ha19f027ca98851ac;
    assign coff[3196] = 64'h5e60fd84a98851ac;
    assign coff[3197] = 64'h05981c26801f4f4f;
    assign coff[3198] = 64'ha98851aca19f027c;
    assign coff[3199] = 64'h801f4f4ffa67e3da;
    assign coff[3200] = 64'h5d2d189aa83ce06e;
    assign coff[3201] = 64'h03d407df800ea8a3;
    assign coff[3202] = 64'ha83ce06ea2d2e766;
    assign coff[3203] = 64'h800ea8a3fc2bf821;
    assign coff[3204] = 64'h7ff1575dfc2bf821;
    assign coff[3205] = 64'h57c31f92a2d2e766;
    assign coff[3206] = 64'hfc2bf821800ea8a3;
    assign coff[3207] = 64'ha2d2e766a83ce06e;
    assign coff[3208] = 64'h77ab2ee2d29344f0;
    assign coff[3209] = 64'h347f97668b42e661;
    assign coff[3210] = 64'hd29344f08854d11e;
    assign coff[3211] = 64'h8b42e661cb80689a;
    assign coff[3212] = 64'h74bd199fcb80689a;
    assign coff[3213] = 64'h2d6cbb108854d11e;
    assign coff[3214] = 64'hcb80689a8b42e661;
    assign coff[3215] = 64'h8854d11ed29344f0;
    assign coff[3216] = 64'h6c81e245bc1a1598;
    assign coff[3217] = 64'h1cb70f4383433314;
    assign coff[3218] = 64'hbc1a1598937e1dbb;
    assign coff[3219] = 64'h83433314e348f0bd;
    assign coff[3220] = 64'h7cbcccece348f0bd;
    assign coff[3221] = 64'h43e5ea68937e1dbb;
    assign coff[3222] = 64'he348f0bd83433314;
    assign coff[3223] = 64'h937e1dbbbc1a1598;
    assign coff[3224] = 64'h7e3b3083eacb56ff;
    assign coff[3225] = 64'h4a43a5b097bf1165;
    assign coff[3226] = 64'heacb56ff81c4cf7d;
    assign coff[3227] = 64'h97bf1165b5bc5a50;
    assign coff[3228] = 64'h6840ee9bb5bc5a50;
    assign coff[3229] = 64'h1534a90181c4cf7d;
    assign coff[3230] = 64'hb5bc5a5097bf1165;
    assign coff[3231] = 64'h81c4cf7deacb56ff;
    assign coff[3232] = 64'h6554666db1cb1304;
    assign coff[3233] = 64'h1059b352810c6f52;
    assign coff[3234] = 64'hb1cb13049aab9993;
    assign coff[3235] = 64'h810c6f52efa64cae;
    assign coff[3236] = 64'h7ef390aeefa64cae;
    assign coff[3237] = 64'h4e34ecfc9aab9993;
    assign coff[3238] = 64'hefa64cae810c6f52;
    assign coff[3239] = 64'h9aab9993b1cb1304;
    assign coff[3240] = 64'h7b8b7b36de8609b1;
    assign coff[3241] = 64'h3fb020ce90f81d7b;
    assign coff[3242] = 64'hde8609b1847484ca;
    assign coff[3243] = 64'h90f81d7bc04fdf32;
    assign coff[3244] = 64'h6f07e285c04fdf32;
    assign coff[3245] = 64'h2179f64f847484ca;
    assign coff[3246] = 64'hc04fdf3290f81d7b;
    assign coff[3247] = 64'h847484cade8609b1;
    assign coff[3248] = 64'h72a3d9f7c7107de4;
    assign coff[3249] = 64'h28cd9fc186ad7e99;
    assign coff[3250] = 64'hc7107de48d5c2609;
    assign coff[3251] = 64'h86ad7e99d732603f;
    assign coff[3252] = 64'h79528167d732603f;
    assign coff[3253] = 64'h38ef821c8d5c2609;
    assign coff[3254] = 64'hd732603f86ad7e99;
    assign coff[3255] = 64'h8d5c2609c7107de4;
    assign coff[3256] = 64'h7fb3af4ef744ec3b;
    assign coff[3257] = 64'h542012e19f870cbc;
    assign coff[3258] = 64'hf744ec3b804c50b2;
    assign coff[3259] = 64'h9f870cbcabdfed1f;
    assign coff[3260] = 64'h6078f344abdfed1f;
    assign coff[3261] = 64'h08bb13c5804c50b2;
    assign coff[3262] = 64'habdfed1f9f870cbc;
    assign coff[3263] = 64'h804c50b2f744ec3b;
    assign coff[3264] = 64'h615ec603acea5af2;
    assign coff[3265] = 64'h0a19fb048066330c;
    assign coff[3266] = 64'hacea5af29ea139fd;
    assign coff[3267] = 64'h8066330cf5e604fc;
    assign coff[3268] = 64'h7f99ccf4f5e604fc;
    assign coff[3269] = 64'h5315a50e9ea139fd;
    assign coff[3270] = 64'hf5e604fc8066330c;
    assign coff[3271] = 64'h9ea139fdacea5af2;
    assign coff[3272] = 64'h79c0e062d880794b;
    assign coff[3273] = 64'h3a29cb918dfa58ea;
    assign coff[3274] = 64'hd880794b863f1f9e;
    assign coff[3275] = 64'h8dfa58eac5d6346f;
    assign coff[3276] = 64'h7205a716c5d6346f;
    assign coff[3277] = 64'h277f86b5863f1f9e;
    assign coff[3278] = 64'hc5d6346f8dfa58ea;
    assign coff[3279] = 64'h863f1f9ed880794b;
    assign coff[3280] = 64'h6fb5507ac182048d;
    assign coff[3281] = 64'h22cd12bd84d25d06;
    assign coff[3282] = 64'hc182048d904aaf86;
    assign coff[3283] = 64'h84d25d06dd32ed43;
    assign coff[3284] = 64'h7b2da2fadd32ed43;
    assign coff[3285] = 64'h3e7dfb73904aaf86;
    assign coff[3286] = 64'hdd32ed4384d25d06;
    assign coff[3287] = 64'h904aaf86c182048d;
    assign coff[3288] = 64'h7f1ea2dcf1038295;
    assign coff[3289] = 64'h4f4a4f899b8412c1;
    assign coff[3290] = 64'hf103829580e15d24;
    assign coff[3291] = 64'h9b8412c1b0b5b077;
    assign coff[3292] = 64'h647bed3fb0b5b077;
    assign coff[3293] = 64'h0efc7d6b80e15d24;
    assign coff[3294] = 64'hb0b5b0779b8412c1;
    assign coff[3295] = 64'h80e15d24f1038295;
    assign coff[3296] = 64'h690b88b5b6dc0685;
    assign coff[3297] = 64'h168f56328200f6ef;
    assign coff[3298] = 64'hb6dc068596f4774b;
    assign coff[3299] = 64'h8200f6efe970a9ce;
    assign coff[3300] = 64'h7dff0911e970a9ce;
    assign coff[3301] = 64'h4923f97b96f4774b;
    assign coff[3302] = 64'he970a9ce8200f6ef;
    assign coff[3303] = 64'h96f4774bb6dc0685;
    assign coff[3304] = 64'h7d09e489e4a03f69;
    assign coff[3305] = 64'h450f2edb943a5bcf;
    assign coff[3306] = 64'he4a03f6982f61b77;
    assign coff[3307] = 64'h943a5bcfbaf0d125;
    assign coff[3308] = 64'h6bc5a431baf0d125;
    assign coff[3309] = 64'h1b5fc09782f61b77;
    assign coff[3310] = 64'hbaf0d125943a5bcf;
    assign coff[3311] = 64'h82f61b77e4a03f69;
    assign coff[3312] = 64'h754bafdcccc21455;
    assign coff[3313] = 64'h2eb502ae88d372c6;
    assign coff[3314] = 64'hccc214558ab45024;
    assign coff[3315] = 64'h88d372c6d14afd52;
    assign coff[3316] = 64'h772c8d3ad14afd52;
    assign coff[3317] = 64'h333debab8ab45024;
    assign coff[3318] = 64'hd14afd5288d372c6;
    assign coff[3319] = 64'h8ab45024ccc21455;
    assign coff[3320] = 64'h7ff9f9ecfd8bb850;
    assign coff[3321] = 64'h58c1f45ba3c585fb;
    assign coff[3322] = 64'hfd8bb85080060614;
    assign coff[3323] = 64'ha3c585fba73e0ba5;
    assign coff[3324] = 64'h5c3a7a05a73e0ba5;
    assign coff[3325] = 64'h027447b080060614;
    assign coff[3326] = 64'ha73e0ba5a3c585fb;
    assign coff[3327] = 64'h80060614fd8bb850;
    assign coff[3328] = 64'h5c179806a719daae;
    assign coff[3329] = 64'h024205e880051939;
    assign coff[3330] = 64'ha719daaea3e867fa;
    assign coff[3331] = 64'h80051939fdbdfa18;
    assign coff[3332] = 64'h7ffae6c7fdbdfa18;
    assign coff[3333] = 64'h58e62552a3e867fa;
    assign coff[3334] = 64'hfdbdfa1880051939;
    assign coff[3335] = 64'ha3e867faa719daae;
    assign coff[3336] = 64'h771a2c88d11c343f;
    assign coff[3337] = 64'h330fd7e18aa039cb;
    assign coff[3338] = 64'hd11c343f88e5d378;
    assign coff[3339] = 64'h8aa039cbccf0281f;
    assign coff[3340] = 64'h755fc635ccf0281f;
    assign coff[3341] = 64'h2ee3cbc188e5d378;
    assign coff[3342] = 64'hccf0281f8aa039cb;
    assign coff[3343] = 64'h88e5d378d11c343f;
    assign coff[3344] = 64'h6baa7d49bac6840c;
    assign coff[3345] = 64'h1b2ea43a82eb652b;
    assign coff[3346] = 64'hbac6840c945582b7;
    assign coff[3347] = 64'h82eb652be4d15bc6;
    assign coff[3348] = 64'h7d149ad5e4d15bc6;
    assign coff[3349] = 64'h45397bf4945582b7;
    assign coff[3350] = 64'he4d15bc682eb652b;
    assign coff[3351] = 64'h945582b7bac6840c;
    assign coff[3352] = 64'h7df62362e93f3107;
    assign coff[3353] = 64'h48fab39196d7c682;
    assign coff[3354] = 64'he93f31078209dc9e;
    assign coff[3355] = 64'h96d7c682b7054c6f;
    assign coff[3356] = 64'h6928397eb7054c6f;
    assign coff[3357] = 64'h16c0cef98209dc9e;
    assign coff[3358] = 64'hb7054c6f96d7c682;
    assign coff[3359] = 64'h8209dc9ee93f3107;
    assign coff[3360] = 64'h645cc260b08e40d2;
    assign coff[3361] = 64'h0eca90ce80db845b;
    assign coff[3362] = 64'hb08e40d29ba33da0;
    assign coff[3363] = 64'h80db845bf1356f32;
    assign coff[3364] = 64'h7f247ba5f1356f32;
    assign coff[3365] = 64'h4f71bf2e9ba33da0;
    assign coff[3366] = 64'hf1356f3280db845b;
    assign coff[3367] = 64'h9ba33da0b08e40d2;
    assign coff[3368] = 64'h7b1feee5dd0290b8;
    assign coff[3369] = 64'h3e52187f90322dbf;
    assign coff[3370] = 64'hdd0290b884e0111b;
    assign coff[3371] = 64'h90322dbfc1ade781;
    assign coff[3372] = 64'h6fcdd241c1ade781;
    assign coff[3373] = 64'h22fd6f4884e0111b;
    assign coff[3374] = 64'hc1ade78190322dbf;
    assign coff[3375] = 64'h84e0111bdd0290b8;
    assign coff[3376] = 64'h71eec716c5a9722c;
    assign coff[3377] = 64'h274fb3ae862fa638;
    assign coff[3378] = 64'hc5a9722c8e1138ea;
    assign coff[3379] = 64'h862fa638d8b04c52;
    assign coff[3380] = 64'h79d059c8d8b04c52;
    assign coff[3381] = 64'h3a568dd48e1138ea;
    assign coff[3382] = 64'hd8b04c52862fa638;
    assign coff[3383] = 64'h8e1138eac5a9722c;
    assign coff[3384] = 64'h7f95cb9af5b3e9f0;
    assign coff[3385] = 64'h52ef61ee9e80a0ee;
    assign coff[3386] = 64'hf5b3e9f0806a3466;
    assign coff[3387] = 64'h9e80a0eead109e12;
    assign coff[3388] = 64'h617f5f12ad109e12;
    assign coff[3389] = 64'h0a4c1610806a3466;
    assign coff[3390] = 64'had109e129e80a0ee;
    assign coff[3391] = 64'h806a3466f5b3e9f0;
    assign coff[3392] = 64'h6057e2a2abba1125;
    assign coff[3393] = 64'h0888ed1b8048ecd5;
    assign coff[3394] = 64'habba11259fa81d5e;
    assign coff[3395] = 64'h8048ecd5f77712e5;
    assign coff[3396] = 64'h7fb7132bf77712e5;
    assign coff[3397] = 64'h5445eedb9fa81d5e;
    assign coff[3398] = 64'hf77712e58048ecd5;
    assign coff[3399] = 64'h9fa81d5eabba1125;
    assign coff[3400] = 64'h79427210d702bec0;
    assign coff[3401] = 64'h38c278d98d45d316;
    assign coff[3402] = 64'hd702bec086bd8df0;
    assign coff[3403] = 64'h8d45d316c73d8727;
    assign coff[3404] = 64'h72ba2ceac73d8727;
    assign coff[3405] = 64'h28fd414086bd8df0;
    assign coff[3406] = 64'hc73d87278d45d316;
    assign coff[3407] = 64'h86bd8df0d702bec0;
    assign coff[3408] = 64'h6eeed758c0244a14;
    assign coff[3409] = 64'h21496fa7846768e7;
    assign coff[3410] = 64'hc0244a14911128a8;
    assign coff[3411] = 64'h846768e7deb69059;
    assign coff[3412] = 64'h7b989719deb69059;
    assign coff[3413] = 64'h3fdbb5ec911128a8;
    assign coff[3414] = 64'hdeb69059846768e7;
    assign coff[3415] = 64'h911128a8c0244a14;
    assign coff[3416] = 64'h7eed1b2cef747365;
    assign coff[3417] = 64'h4e0d1c309a8ceb31;
    assign coff[3418] = 64'hef7473658112e4d4;
    assign coff[3419] = 64'h9a8ceb31b1f2e3d0;
    assign coff[3420] = 64'h657314cfb1f2e3d0;
    assign coff[3421] = 64'h108b8c9b8112e4d4;
    assign coff[3422] = 64'hb1f2e3d09a8ceb31;
    assign coff[3423] = 64'h8112e4d4ef747365;
    assign coff[3424] = 64'h6823bcb7b5936f53;
    assign coff[3425] = 64'h1503153a81bc8564;
    assign coff[3426] = 64'hb5936f5397dc4349;
    assign coff[3427] = 64'h81bc8564eafceac6;
    assign coff[3428] = 64'h7e437a9ceafceac6;
    assign coff[3429] = 64'h4a6c90ad97dc4349;
    assign coff[3430] = 64'heafceac681bc8564;
    assign coff[3431] = 64'h97dc4349b5936f53;
    assign coff[3432] = 64'h7cb17c8de317f6fa;
    assign coff[3433] = 64'h43bb48d493637c3d;
    assign coff[3434] = 64'he317f6fa834e8373;
    assign coff[3435] = 64'h93637c3dbc44b72c;
    assign coff[3436] = 64'h6c9c83c3bc44b72c;
    assign coff[3437] = 64'h1ce80906834e8373;
    assign coff[3438] = 64'hbc44b72c93637c3d;
    assign coff[3439] = 64'h834e8373e317f6fa;
    assign coff[3440] = 64'h74a872e8cb5294ce;
    assign coff[3441] = 64'h2d3db928884303c1;
    assign coff[3442] = 64'hcb5294ce8b578d18;
    assign coff[3443] = 64'h884303c1d2c246d8;
    assign coff[3444] = 64'h77bcfc3fd2c246d8;
    assign coff[3445] = 64'h34ad6b328b578d18;
    assign coff[3446] = 64'hd2c246d8884303c1;
    assign coff[3447] = 64'h8b578d18cb5294ce;
    assign coff[3448] = 64'h7fefcca4fbf9ba39;
    assign coff[3449] = 64'h579e81b8a2b077c5;
    assign coff[3450] = 64'hfbf9ba398010335c;
    assign coff[3451] = 64'ha2b077c5a8617e48;
    assign coff[3452] = 64'h5d4f883ba8617e48;
    assign coff[3453] = 64'h040645c78010335c;
    assign coff[3454] = 64'ha8617e48a2b077c5;
    assign coff[3455] = 64'h8010335cfbf9ba39;
    assign coff[3456] = 64'h5e3f0194a9634858;
    assign coff[3457] = 64'h0565e40d801d26c8;
    assign coff[3458] = 64'ha9634858a1c0fe6c;
    assign coff[3459] = 64'h801d26c8fa9a1bf3;
    assign coff[3460] = 64'h7fe2d938fa9a1bf3;
    assign coff[3461] = 64'h569cb7a8a1c0fe6c;
    assign coff[3462] = 64'hfa9a1bf3801d26c8;
    assign coff[3463] = 64'ha1c0fe6ca9634858;
    assign coff[3464] = 64'h7837942bd40c15f3;
    assign coff[3465] = 64'h35ed50c98bea131e;
    assign coff[3466] = 64'hd40c15f387c86bd5;
    assign coff[3467] = 64'h8bea131eca12af37;
    assign coff[3468] = 64'h7415ece2ca12af37;
    assign coff[3469] = 64'h2bf3ea0d87c86bd5;
    assign coff[3470] = 64'hca12af378bea131e;
    assign coff[3471] = 64'h87c86bd5d40c15f3;
    assign coff[3472] = 64'h6d551858bd704542;
    assign coff[3473] = 64'h1e3e5ee5839fd014;
    assign coff[3474] = 64'hbd70454292aae7a8;
    assign coff[3475] = 64'h839fd014e1c1a11b;
    assign coff[3476] = 64'h7c602fece1c1a11b;
    assign coff[3477] = 64'h428fbabe92aae7a8;
    assign coff[3478] = 64'he1c1a11b839fd014;
    assign coff[3479] = 64'h92aae7a8bd704542;
    assign coff[3480] = 64'h7e7b5fceec584e41;
    assign coff[3481] = 64'h4b89badd98aa6136;
    assign coff[3482] = 64'hec584e418184a032;
    assign coff[3483] = 64'h98aa6136b4764523;
    assign coff[3484] = 64'h67559ecab4764523;
    assign coff[3485] = 64'h13a7b1bf8184a032;
    assign coff[3486] = 64'hb476452398aa6136;
    assign coff[3487] = 64'h8184a032ec584e41;
    assign coff[3488] = 64'h66482267b30ae912;
    assign coff[3489] = 64'h11e8347881423f3a;
    assign coff[3490] = 64'hb30ae91299b7dd99;
    assign coff[3491] = 64'h81423f3aee17cb88;
    assign coff[3492] = 64'h7ebdc0c6ee17cb88;
    assign coff[3493] = 64'h4cf516ee99b7dd99;
    assign coff[3494] = 64'hee17cb8881423f3a;
    assign coff[3495] = 64'h99b7dd99b30ae912;
    assign coff[3496] = 64'h7bf24434e00acd0e;
    assign coff[3497] = 64'h410bb48c91c25508;
    assign coff[3498] = 64'he00acd0e840dbbcc;
    assign coff[3499] = 64'h91c25508bef44b74;
    assign coff[3500] = 64'h6e3daaf8bef44b74;
    assign coff[3501] = 64'h1ff532f2840dbbcc;
    assign coff[3502] = 64'hbef44b7491c25508;
    assign coff[3503] = 64'h840dbbcce00acd0e;
    assign coff[3504] = 64'h73548168c879bb89;
    assign coff[3505] = 64'h2a49f9208730045d;
    assign coff[3506] = 64'hc879bb898cab7e98;
    assign coff[3507] = 64'h8730045dd5b606e0;
    assign coff[3508] = 64'h78cffba3d5b606e0;
    assign coff[3509] = 64'h378644778cab7e98;
    assign coff[3510] = 64'hd5b606e08730045d;
    assign coff[3511] = 64'h8cab7e98c879bb89;
    assign coff[3512] = 64'h7fcca6a7f8d644b2;
    assign coff[3513] = 64'h554d858da09130ad;
    assign coff[3514] = 64'hf8d644b280335959;
    assign coff[3515] = 64'ha09130adaab27a73;
    assign coff[3516] = 64'h5f6ecf53aab27a73;
    assign coff[3517] = 64'h0729bb4e80335959;
    assign coff[3518] = 64'haab27a73a09130ad;
    assign coff[3519] = 64'h80335959f8d644b2;
    assign coff[3520] = 64'h6261e866ae1dd8c0;
    assign coff[3521] = 64'h0baaa53b8088649e;
    assign coff[3522] = 64'hae1dd8c09d9e179a;
    assign coff[3523] = 64'h8088649ef4555ac5;
    assign coff[3524] = 64'h7f779b62f4555ac5;
    assign coff[3525] = 64'h51e227409d9e179a;
    assign coff[3526] = 64'hf4555ac58088649e;
    assign coff[3527] = 64'h9d9e179aae1dd8c0;
    assign coff[3528] = 64'h7a3a9d0fd9ffb9a9;
    assign coff[3529] = 64'h3b8ee03e8eb34415;
    assign coff[3530] = 64'hd9ffb9a985c562f1;
    assign coff[3531] = 64'h8eb34415c4711fc2;
    assign coff[3532] = 64'h714cbbebc4711fc2;
    assign coff[3533] = 64'h2600465785c562f1;
    assign coff[3534] = 64'hc4711fc28eb34415;
    assign coff[3535] = 64'h85c562f1d9ffb9a9;
    assign coff[3536] = 64'h70777b1cc2e227cb;
    assign coff[3537] = 64'h244f5e5c854210db;
    assign coff[3538] = 64'hc2e227cb8f8884e4;
    assign coff[3539] = 64'h854210dbdbb0a1a4;
    assign coff[3540] = 64'h7abdef25dbb0a1a4;
    assign coff[3541] = 64'h3d1dd8358f8884e4;
    assign coff[3542] = 64'hdbb0a1a4854210db;
    assign coff[3543] = 64'h8f8884e4c2e227cb;
    assign coff[3544] = 64'h7f4b43f2f29325ad;
    assign coff[3545] = 64'h508474549c7f1a0a;
    assign coff[3546] = 64'hf29325ad80b4bc0e;
    assign coff[3547] = 64'h9c7f1a0aaf7b8bac;
    assign coff[3548] = 64'h6380e5f6af7b8bac;
    assign coff[3549] = 64'h0d6cda5380b4bc0e;
    assign coff[3550] = 64'haf7b8bac9c7f1a0a;
    assign coff[3551] = 64'h80b4bc0ef29325ad;
    assign coff[3552] = 64'h69ef47f6b8276f93;
    assign coff[3553] = 64'h181ab881824a43fe;
    assign coff[3554] = 64'hb8276f939610b80a;
    assign coff[3555] = 64'h824a43fee7e5477f;
    assign coff[3556] = 64'h7db5bc02e7e5477f;
    assign coff[3557] = 64'h47d8906d9610b80a;
    assign coff[3558] = 64'he7e5477f824a43fe;
    assign coff[3559] = 64'h9610b80ab8276f93;
    assign coff[3560] = 64'h7d5d7a74e6299604;
    assign coff[3561] = 64'h46606b4e95156308;
    assign coff[3562] = 64'he629960482a2858c;
    assign coff[3563] = 64'h95156308b99f94b2;
    assign coff[3564] = 64'h6aea9cf8b99f94b2;
    assign coff[3565] = 64'h19d669fc82a2858c;
    assign coff[3566] = 64'hb99f94b295156308;
    assign coff[3567] = 64'h82a2858ce6299604;
    assign coff[3568] = 64'h75ea672ace338d97;
    assign coff[3569] = 64'h302a7f3a896879fb;
    assign coff[3570] = 64'hce338d978a1598d6;
    assign coff[3571] = 64'h896879fbcfd580c6;
    assign coff[3572] = 64'h76978605cfd580c6;
    assign coff[3573] = 64'h31cc72698a1598d6;
    assign coff[3574] = 64'hcfd580c6896879fb;
    assign coff[3575] = 64'h8a1598d6ce338d97;
    assign coff[3576] = 64'h7fff3824ff1dcea0;
    assign coff[3577] = 64'h59e1faffa4de2270;
    assign coff[3578] = 64'hff1dcea08000c7dc;
    assign coff[3579] = 64'ha4de2270a61e0501;
    assign coff[3580] = 64'h5b21dd90a61e0501;
    assign coff[3581] = 64'h00e231608000c7dc;
    assign coff[3582] = 64'ha61e0501a4de2270;
    assign coff[3583] = 64'h8000c7dcff1dcea0;
    assign coff[3584] = 64'h5b8b8239a689a022;
    assign coff[3585] = 64'h0178fb9980022b29;
    assign coff[3586] = 64'ha689a022a4747dc7;
    assign coff[3587] = 64'h80022b29fe870467;
    assign coff[3588] = 64'h7ffdd4d7fe870467;
    assign coff[3589] = 64'h59765fdea4747dc7;
    assign coff[3590] = 64'hfe87046780022b29;
    assign coff[3591] = 64'ha4747dc7a689a022;
    assign coff[3592] = 64'h76cff232d061588b;
    assign coff[3593] = 64'h32573a3f8a509585;
    assign coff[3594] = 64'hd061588b89300dce;
    assign coff[3595] = 64'h8a509585cda8c5c1;
    assign coff[3596] = 64'h75af6a7bcda8c5c1;
    assign coff[3597] = 64'h2f9ea77589300dce;
    assign coff[3598] = 64'hcda8c5c18a509585;
    assign coff[3599] = 64'h89300dced061588b;
    assign coff[3600] = 64'h6b3d3bcbba1dbaaa;
    assign coff[3601] = 64'h1a6a092982c14cf1;
    assign coff[3602] = 64'hba1dbaaa94c2c435;
    assign coff[3603] = 64'h82c14cf1e595f6d7;
    assign coff[3604] = 64'h7d3eb30fe595f6d7;
    assign coff[3605] = 64'h45e2455694c2c435;
    assign coff[3606] = 64'he595f6d782c14cf1;
    assign coff[3607] = 64'h94c2c435ba1dbaaa;
    assign coff[3608] = 64'h7dd1ca75e879714d;
    assign coff[3609] = 64'h48552b9b9665a5b4;
    assign coff[3610] = 64'he879714d822e358b;
    assign coff[3611] = 64'h9665a5b4b7aad465;
    assign coff[3612] = 64'h699a5a4cb7aad465;
    assign coff[3613] = 64'h17868eb3822e358b;
    assign coff[3614] = 64'hb7aad4659665a5b4;
    assign coff[3615] = 64'h822e358be879714d;
    assign coff[3616] = 64'h63df7c4daff0fcfe;
    assign coff[3617] = 64'h0e02c7d780c4e553;
    assign coff[3618] = 64'haff0fcfe9c2083b3;
    assign coff[3619] = 64'h80c4e553f1fd3829;
    assign coff[3620] = 64'h7f3b1aadf1fd3829;
    assign coff[3621] = 64'h500f03029c2083b3;
    assign coff[3622] = 64'hf1fd382980c4e553;
    assign coff[3623] = 64'h9c2083b3aff0fcfe;
    assign coff[3624] = 64'h7ae860c7dc4154cd;
    assign coff[3625] = 64'h3da22cd78fd0d333;
    assign coff[3626] = 64'hdc4154cd85179f39;
    assign coff[3627] = 64'h8fd0d333c25dd329;
    assign coff[3628] = 64'h702f2ccdc25dd329;
    assign coff[3629] = 64'h23beab3385179f39;
    assign coff[3630] = 64'hc25dd3298fd0d333;
    assign coff[3631] = 64'h85179f39dc4154cd;
    assign coff[3632] = 64'h71929789c4f6c35d;
    assign coff[3633] = 64'h26902b3985f27c93;
    assign coff[3634] = 64'hc4f6c35d8e6d6877;
    assign coff[3635] = 64'h85f27c93d96fd4c7;
    assign coff[3636] = 64'h7a0d836dd96fd4c7;
    assign coff[3637] = 64'h3b093ca38e6d6877;
    assign coff[3638] = 64'hd96fd4c785f27c93;
    assign coff[3639] = 64'h8e6d6877c4f6c35d;
    assign coff[3640] = 64'h7f850179f4eb8def;
    assign coff[3641] = 64'h5255d5c59dfed33e;
    assign coff[3642] = 64'hf4eb8def807afe87;
    assign coff[3643] = 64'h9dfed33eadaa2a3b;
    assign coff[3644] = 64'h62012cc2adaa2a3b;
    assign coff[3645] = 64'h0b147211807afe87;
    assign coff[3646] = 64'hadaa2a3b9dfed33e;
    assign coff[3647] = 64'h807afe87f4eb8def;
    assign coff[3648] = 64'h5fd30bbcab23236a;
    assign coff[3649] = 64'h07c04598803c2257;
    assign coff[3650] = 64'hab23236aa02cf444;
    assign coff[3651] = 64'h803c2257f83fba68;
    assign coff[3652] = 64'h7fc3dda9f83fba68;
    assign coff[3653] = 64'h54dcdc96a02cf444;
    assign coff[3654] = 64'hf83fba68803c2257;
    assign coff[3655] = 64'ha02cf444ab23236a;
    assign coff[3656] = 64'h790179cdd6447844;
    assign coff[3657] = 64'h380dfc8d8ced385b;
    assign coff[3658] = 64'hd644784486fe8633;
    assign coff[3659] = 64'h8ced385bc7f20373;
    assign coff[3660] = 64'h7312c7a5c7f20373;
    assign coff[3661] = 64'h29bb87bc86fe8633;
    assign coff[3662] = 64'hc7f203738ced385b;
    assign coff[3663] = 64'h86fe8633d6447844;
    assign coff[3664] = 64'h6e89ffb9bf765858;
    assign coff[3665] = 64'h208721f98433b806;
    assign coff[3666] = 64'hbf76585891760047;
    assign coff[3667] = 64'h8433b806df78de07;
    assign coff[3668] = 64'h7bcc47fadf78de07;
    assign coff[3669] = 64'h4089a7a891760047;
    assign coff[3670] = 64'hdf78de078433b806;
    assign coff[3671] = 64'h91760047bf765858;
    assign coff[3672] = 64'h7ed28171eead2813;
    assign coff[3673] = 64'h4d6d60df9a12ce4b;
    assign coff[3674] = 64'heead2813812d7e8f;
    assign coff[3675] = 64'h9a12ce4bb2929f21;
    assign coff[3676] = 64'h65ed31b5b2929f21;
    assign coff[3677] = 64'h1152d7ed812d7e8f;
    assign coff[3678] = 64'hb2929f219a12ce4b;
    assign coff[3679] = 64'h812d7e8feead2813;
    assign coff[3680] = 64'h67ae54bab4f03663;
    assign coff[3681] = 64'h143ca605819c1fc5;
    assign coff[3682] = 64'hb4f036639851ab46;
    assign coff[3683] = 64'h819c1fc5ebc359fb;
    assign coff[3684] = 64'h7e63e03bebc359fb;
    assign coff[3685] = 64'h4b0fc99d9851ab46;
    assign coff[3686] = 64'hebc359fb819c1fc5;
    assign coff[3687] = 64'h9851ab46b4f03663;
    assign coff[3688] = 64'h7c837ad8e2543ccc;
    assign coff[3689] = 64'h43105a5092f99deb;
    assign coff[3690] = 64'he2543ccc837c8528;
    assign coff[3691] = 64'h92f99debbcefa5b0;
    assign coff[3692] = 64'h6d066215bcefa5b0;
    assign coff[3693] = 64'h1dabc334837c8528;
    assign coff[3694] = 64'hbcefa5b092f99deb;
    assign coff[3695] = 64'h837c8528e2543ccc;
    assign coff[3696] = 64'h74552446ca9b971e;
    assign coff[3697] = 64'h2c816c0c87fc870f;
    assign coff[3698] = 64'hca9b971e8baadbba;
    assign coff[3699] = 64'h87fc870fd37e93f4;
    assign coff[3700] = 64'h780378f1d37e93f4;
    assign coff[3701] = 64'h356468e28baadbba;
    assign coff[3702] = 64'hd37e93f487fc870f;
    assign coff[3703] = 64'h8baadbbaca9b971e;
    assign coff[3704] = 64'h7fe8dc78fb30c91b;
    assign coff[3705] = 64'h570b8369a2274959;
    assign coff[3706] = 64'hfb30c91b80172388;
    assign coff[3707] = 64'ha2274959a8f47c97;
    assign coff[3708] = 64'h5dd8b6a7a8f47c97;
    assign coff[3709] = 64'h04cf36e580172388;
    assign coff[3710] = 64'ha8f47c97a2274959;
    assign coff[3711] = 64'h80172388fb30c91b;
    assign coff[3712] = 64'h5db680b4a8cfa8d2;
    assign coff[3713] = 64'h049cfba7801549e6;
    assign coff[3714] = 64'ha8cfa8d2a2497f4c;
    assign coff[3715] = 64'h801549e6fb630459;
    assign coff[3716] = 64'h7feab61afb630459;
    assign coff[3717] = 64'h5730572ea2497f4c;
    assign coff[3718] = 64'hfb630459801549e6;
    assign coff[3719] = 64'ha2497f4ca8cfa8d2;
    assign coff[3720] = 64'h77f1f581d34f764f;
    assign coff[3721] = 64'h3536b5be8b95ed21;
    assign coff[3722] = 64'hd34f764f880e0a7f;
    assign coff[3723] = 64'h8b95ed21cac94a42;
    assign coff[3724] = 64'h746a12dfcac94a42;
    assign coff[3725] = 64'h2cb089b1880e0a7f;
    assign coff[3726] = 64'hcac94a428b95ed21;
    assign coff[3727] = 64'h880e0a7fd34f764f;
    assign coff[3728] = 64'h6cec03afbcc4da7b;
    assign coff[3729] = 64'h1d7adb738370e7e9;
    assign coff[3730] = 64'hbcc4da7b9313fc51;
    assign coff[3731] = 64'h8370e7e9e285248d;
    assign coff[3732] = 64'h7c8f1817e285248d;
    assign coff[3733] = 64'h433b25859313fc51;
    assign coff[3734] = 64'he285248d8370e7e9;
    assign coff[3735] = 64'h9313fc51bcc4da7b;
    assign coff[3736] = 64'h7e5be40ceb91b96c;
    assign coff[3737] = 64'h4ae70caf98343940;
    assign coff[3738] = 64'heb91b96c81a41bf4;
    assign coff[3739] = 64'h98343940b518f351;
    assign coff[3740] = 64'h67cbc6c0b518f351;
    assign coff[3741] = 64'h146e469481a41bf4;
    assign coff[3742] = 64'hb518f35198343940;
    assign coff[3743] = 64'h81a41bf4eb91b96c;
    assign coff[3744] = 64'h65cec204b26a9e54;
    assign coff[3745] = 64'h112109078126bac8;
    assign coff[3746] = 64'hb26a9e549a313dfc;
    assign coff[3747] = 64'h8126bac8eedef6f9;
    assign coff[3748] = 64'h7ed94538eedef6f9;
    assign coff[3749] = 64'h4d9561ac9a313dfc;
    assign coff[3750] = 64'heedef6f98126bac8;
    assign coff[3751] = 64'h9a313dfcb26a9e54;
    assign coff[3752] = 64'h7bbf7860df484302;
    assign coff[3753] = 64'h405e3a16915cb0c3;
    assign coff[3754] = 64'hdf484302844087a0;
    assign coff[3755] = 64'h915cb0c3bfa1c5ea;
    assign coff[3756] = 64'h6ea34f3dbfa1c5ea;
    assign coff[3757] = 64'h20b7bcfe844087a0;
    assign coff[3758] = 64'hbfa1c5ea915cb0c3;
    assign coff[3759] = 64'h844087a0df484302;
    assign coff[3760] = 64'h72fcbb8cc7c4d757;
    assign coff[3761] = 64'h298bffb286ee2c1e;
    assign coff[3762] = 64'hc7c4d7578d034474;
    assign coff[3763] = 64'h86ee2c1ed674004e;
    assign coff[3764] = 64'h7911d3e2d674004e;
    assign coff[3765] = 64'h383b28a98d034474;
    assign coff[3766] = 64'hd674004e86ee2c1e;
    assign coff[3767] = 64'h8d034474c7c4d757;
    assign coff[3768] = 64'h7fc0c896f80d8ea9;
    assign coff[3769] = 64'h54b734baa00ba853;
    assign coff[3770] = 64'hf80d8ea9803f376a;
    assign coff[3771] = 64'ha00ba853ab48cb46;
    assign coff[3772] = 64'h5ff457adab48cb46;
    assign coff[3773] = 64'h07f27157803f376a;
    assign coff[3774] = 64'hab48cb46a00ba853;
    assign coff[3775] = 64'h803f376af80d8ea9;
    assign coff[3776] = 64'h61e0cff5ad83b416;
    assign coff[3777] = 64'h0ae25d8d8076ae7e;
    assign coff[3778] = 64'had83b4169e1f300b;
    assign coff[3779] = 64'h8076ae7ef51da273;
    assign coff[3780] = 64'h7f895182f51da273;
    assign coff[3781] = 64'h527c4bea9e1f300b;
    assign coff[3782] = 64'hf51da2738076ae7e;
    assign coff[3783] = 64'h9e1f300bad83b416;
    assign coff[3784] = 64'h79fe5539d93fe9ab;
    assign coff[3785] = 64'h3adc9e868e564246;
    assign coff[3786] = 64'hd93fe9ab8601aac7;
    assign coff[3787] = 64'h8e564246c523617a;
    assign coff[3788] = 64'h71a9bdbac523617a;
    assign coff[3789] = 64'h26c016558601aac7;
    assign coff[3790] = 64'hc523617a8e564246;
    assign coff[3791] = 64'h8601aac7d93fe9ab;
    assign coff[3792] = 64'h7016f014c231c9ec;
    assign coff[3793] = 64'h238e646a85099f3e;
    assign coff[3794] = 64'hc231c9ec8fe90fec;
    assign coff[3795] = 64'h85099f3edc719b96;
    assign coff[3796] = 64'h7af660c2dc719b96;
    assign coff[3797] = 64'h3dce36148fe90fec;
    assign coff[3798] = 64'hdc719b9685099f3e;
    assign coff[3799] = 64'h8fe90fecc231c9ec;
    assign coff[3800] = 64'h7f359057f1cb429a;
    assign coff[3801] = 64'h4fe7c4839c011b08;
    assign coff[3802] = 64'hf1cb429a80ca6fa9;
    assign coff[3803] = 64'h9c011b08b0183b7d;
    assign coff[3804] = 64'h63fee4f8b0183b7d;
    assign coff[3805] = 64'h0e34bd6680ca6fa9;
    assign coff[3806] = 64'hb0183b7d9c011b08;
    assign coff[3807] = 64'h80ca6fa9f1cb429a;
    assign coff[3808] = 64'h697dea7bb781619c;
    assign coff[3809] = 64'h1755242282250232;
    assign coff[3810] = 64'hb781619c96821585;
    assign coff[3811] = 64'h82250232e8aadbde;
    assign coff[3812] = 64'h7ddafdcee8aadbde;
    assign coff[3813] = 64'h487e9e6496821585;
    assign coff[3814] = 64'he8aadbde82250232;
    assign coff[3815] = 64'h96821585b781619c;
    assign coff[3816] = 64'h7d3449f5e564c9e3;
    assign coff[3817] = 64'h45b8231894a75afd;
    assign coff[3818] = 64'he564c9e382cbb60b;
    assign coff[3819] = 64'h94a75afdba47dce8;
    assign coff[3820] = 64'h6b58a503ba47dce8;
    assign coff[3821] = 64'h1a9b361d82cbb60b;
    assign coff[3822] = 64'hba47dce894a75afd;
    assign coff[3823] = 64'h82cbb60be564c9e3;
    assign coff[3824] = 64'h759b9c9bcd7a92a2;
    assign coff[3825] = 64'h2f6ffb7a891d63b5;
    assign coff[3826] = 64'hcd7a92a28a646365;
    assign coff[3827] = 64'h891d63b5d0900486;
    assign coff[3828] = 64'h76e29c4bd0900486;
    assign coff[3829] = 64'h32856d5e8a646365;
    assign coff[3830] = 64'hd0900486891d63b5;
    assign coff[3831] = 64'h8a646365cd7a92a2;
    assign coff[3832] = 64'h7ffd36eefe54c169;
    assign coff[3833] = 64'h595265dfa4516319;
    assign coff[3834] = 64'hfe54c1698002c912;
    assign coff[3835] = 64'ha4516319a6ad9a21;
    assign coff[3836] = 64'h5bae9ce7a6ad9a21;
    assign coff[3837] = 64'h01ab3e978002c912;
    assign coff[3838] = 64'ha6ad9a21a4516319;
    assign coff[3839] = 64'h8002c912fe54c169;
    assign coff[3840] = 64'h5ca2ca99a7aaf094;
    assign coff[3841] = 64'h030b0aa480094310;
    assign coff[3842] = 64'ha7aaf094a35d3567;
    assign coff[3843] = 64'h80094310fcf4f55c;
    assign coff[3844] = 64'h7ff6bcf0fcf4f55c;
    assign coff[3845] = 64'h58550f6ca35d3567;
    assign coff[3846] = 64'hfcf4f55c80094310;
    assign coff[3847] = 64'ha35d3567a7aaf094;
    assign coff[3848] = 64'h776340ffd1d783a6;
    assign coff[3849] = 64'h33c7f7858af0ffac;
    assign coff[3850] = 64'hd1d783a6889cbf01;
    assign coff[3851] = 64'h8af0ffaccc38087b;
    assign coff[3852] = 64'h750f0054cc38087b;
    assign coff[3853] = 64'h2e287c5a889cbf01;
    assign coff[3854] = 64'hcc38087b8af0ffac;
    assign coff[3855] = 64'h889cbf01d1d783a6;
    assign coff[3856] = 64'h6c16b521bb6ff83c;
    assign coff[3857] = 64'h1bf2fc3a8316b205;
    assign coff[3858] = 64'hbb6ff83c93e94adf;
    assign coff[3859] = 64'h8316b205e40d03c6;
    assign coff[3860] = 64'h7ce94dfbe40d03c6;
    assign coff[3861] = 64'h449007c493e94adf;
    assign coff[3862] = 64'he40d03c68316b205;
    assign coff[3863] = 64'h93e94adfbb6ff83c;
    assign coff[3864] = 64'h7e194584ea0528e5;
    assign coff[3865] = 64'h499f8774974aeac6;
    assign coff[3866] = 64'hea0528e581e6ba7c;
    assign coff[3867] = 64'h974aeac6b660788c;
    assign coff[3868] = 64'h68b5153ab660788c;
    assign coff[3869] = 64'h15fad71b81e6ba7c;
    assign coff[3870] = 64'hb660788c974aeac6;
    assign coff[3871] = 64'h81e6ba7cea0528e5;
    assign coff[3872] = 64'h64d910d1b12c48ab;
    assign coff[3873] = 64'h0f92354680f35d19;
    assign coff[3874] = 64'hb12c48ab9b26ef2f;
    assign coff[3875] = 64'h80f35d19f06dcaba;
    assign coff[3876] = 64'h7f0ca2e7f06dcaba;
    assign coff[3877] = 64'h4ed3b7559b26ef2f;
    assign coff[3878] = 64'hf06dcaba80f35d19;
    assign coff[3879] = 64'h9b26ef2fb12c48ab;
    assign coff[3880] = 64'h7b564d36ddc422f8;
    assign coff[3881] = 64'h3f016a6190949c28;
    assign coff[3882] = 64'hddc422f884a9b2ca;
    assign coff[3883] = 64'h90949c28c0fe959f;
    assign coff[3884] = 64'h6f6b63d8c0fe959f;
    assign coff[3885] = 64'h223bdd0884a9b2ca;
    assign coff[3886] = 64'hc0fe959f90949c28;
    assign coff[3887] = 64'h84a9b2caddc422f8;
    assign coff[3888] = 64'h7249dd86c65cb0ed;
    assign coff[3889] = 64'h280edb23866dfc6e;
    assign coff[3890] = 64'hc65cb0ed8db6227a;
    assign coff[3891] = 64'h866dfc6ed7f124dd;
    assign coff[3892] = 64'h79920392d7f124dd;
    assign coff[3893] = 64'h39a34f138db6227a;
    assign coff[3894] = 64'hd7f124dd866dfc6e;
    assign coff[3895] = 64'h8db6227ac65cb0ed;
    assign coff[3896] = 64'h7fa55aeef67c5f59;
    assign coff[3897] = 64'h538821759f035f2e;
    assign coff[3898] = 64'hf67c5f59805aa512;
    assign coff[3899] = 64'h9f035f2eac77de8b;
    assign coff[3900] = 64'h60fca0d2ac77de8b;
    assign coff[3901] = 64'h0983a0a7805aa512;
    assign coff[3902] = 64'hac77de8b9f035f2e;
    assign coff[3903] = 64'h805aa512f67c5f59;
    assign coff[3904] = 64'h60dbcbd1ac51cecf;
    assign coff[3905] = 64'h09517f8f8056f272;
    assign coff[3906] = 64'hac51cecf9f24342f;
    assign coff[3907] = 64'h8056f272f6ae8071;
    assign coff[3908] = 64'h7fa90d8ef6ae8071;
    assign coff[3909] = 64'h53ae31319f24342f;
    assign coff[3910] = 64'hf6ae80718056f272;
    assign coff[3911] = 64'h9f24342fac51cecf;
    assign coff[3912] = 64'h79823f20d7c16a5f;
    assign coff[3913] = 64'h397669198d9f88e5;
    assign coff[3914] = 64'hd7c16a5f867dc0e0;
    assign coff[3915] = 64'h8d9f88e5c68996e7;
    assign coff[3916] = 64'h7260771bc68996e7;
    assign coff[3917] = 64'h283e95a1867dc0e0;
    assign coff[3918] = 64'hc68996e78d9f88e5;
    assign coff[3919] = 64'h867dc0e0d7c16a5f;
    assign coff[3920] = 64'h6f529d40c0d2d960;
    assign coff[3921] = 64'h220b6b32849c4abd;
    assign coff[3922] = 64'hc0d2d96090ad62c0;
    assign coff[3923] = 64'h849c4abdddf494ce;
    assign coff[3924] = 64'h7b63b543ddf494ce;
    assign coff[3925] = 64'h3f2d26a090ad62c0;
    assign coff[3926] = 64'hddf494ce849c4abd;
    assign coff[3927] = 64'h90ad62c0c0d2d960;
    assign coff[3928] = 64'h7f067bbaf03be78a;
    assign coff[3929] = 64'h4eac16eb9b080268;
    assign coff[3930] = 64'hf03be78a80f98446;
    assign coff[3931] = 64'h9b080268b153e915;
    assign coff[3932] = 64'h64f7fd98b153e915;
    assign coff[3933] = 64'h0fc4187680f98446;
    assign coff[3934] = 64'hb153e9159b080268;
    assign coff[3935] = 64'h80f98446f03be78a;
    assign coff[3936] = 64'h689823bfb6375fe5;
    assign coff[3937] = 64'h15c9509781de228d;
    assign coff[3938] = 64'hb6375fe59767dc41;
    assign coff[3939] = 64'h81de228dea36af69;
    assign coff[3940] = 64'h7e21dd73ea36af69;
    assign coff[3941] = 64'h49c8a01b9767dc41;
    assign coff[3942] = 64'hea36af6981de228d;
    assign coff[3943] = 64'h9767dc41b6375fe5;
    assign coff[3944] = 64'h7cde4a98e3dbf87a;
    assign coff[3945] = 64'h4465903993ce668b;
    assign coff[3946] = 64'he3dbf87a8321b568;
    assign coff[3947] = 64'h93ce668bbb9a6fc7;
    assign coff[3948] = 64'h6c319975bb9a6fc7;
    assign coff[3949] = 64'h1c2407868321b568;
    assign coff[3950] = 64'hbb9a6fc793ce668b;
    assign coff[3951] = 64'h8321b568e3dbf87a;
    assign coff[3952] = 64'h74faa1b3cc0a1477;
    assign coff[3953] = 64'h2df996a3888aa7e3;
    assign coff[3954] = 64'hcc0a14778b055e4d;
    assign coff[3955] = 64'h888aa7e3d206695d;
    assign coff[3956] = 64'h7775581dd206695d;
    assign coff[3957] = 64'h33f5eb898b055e4d;
    assign coff[3958] = 64'hd206695d888aa7e3;
    assign coff[3959] = 64'h8b055e4dcc0a1477;
    assign coff[3960] = 64'h7ff58125fcc2b545;
    assign coff[3961] = 64'h5830a7d6a33a8c6c;
    assign coff[3962] = 64'hfcc2b545800a7edb;
    assign coff[3963] = 64'ha33a8c6ca7cf582a;
    assign coff[3964] = 64'h5cc57394a7cf582a;
    assign coff[3965] = 64'h033d4abb800a7edb;
    assign coff[3966] = 64'ha7cf582aa33a8c6c;
    assign coff[3967] = 64'h800a7edbfcc2b545;
    assign coff[3968] = 64'h5ec699e9a9f7bd92;
    assign coff[3969] = 64'h062ebf2280263f36;
    assign coff[3970] = 64'ha9f7bd92a1396617;
    assign coff[3971] = 64'h80263f36f9d140de;
    assign coff[3972] = 64'h7fd9c0caf9d140de;
    assign coff[3973] = 64'h5608426ea1396617;
    assign coff[3974] = 64'hf9d140de80263f36;
    assign coff[3975] = 64'ha1396617a9f7bd92;
    assign coff[3976] = 64'h787c0a36d4c92209;
    assign coff[3977] = 64'h36a366c68c3f5788;
    assign coff[3978] = 64'hd4c922098783f5ca;
    assign coff[3979] = 64'h8c3f5788c95c993a;
    assign coff[3980] = 64'h73c0a878c95c993a;
    assign coff[3981] = 64'h2b36ddf78783f5ca;
    assign coff[3982] = 64'hc95c993a8c3f5788;
    assign coff[3983] = 64'h8783f5cad4c92209;
    assign coff[3984] = 64'h6dbd1f3cbe1c5444;
    assign coff[3985] = 64'h1f0197b883cfeb22;
    assign coff[3986] = 64'hbe1c54449242e0c4;
    assign coff[3987] = 64'h83cfeb22e0fe6848;
    assign coff[3988] = 64'h7c3014dee0fe6848;
    assign coff[3989] = 64'h41e3abbc9242e0c4;
    assign coff[3990] = 64'he0fe684883cfeb22;
    assign coff[3991] = 64'h9242e0c4be1c5444;
    assign coff[3992] = 64'h7e99a37ced1f1396;
    assign coff[3993] = 64'h4c2baea999218824;
    assign coff[3994] = 64'hed1f139681665c84;
    assign coff[3995] = 64'h99218824b3d45157;
    assign coff[3996] = 64'h66de77dcb3d45157;
    assign coff[3997] = 64'h12e0ec6a81665c84;
    assign coff[3998] = 64'hb3d4515799218824;
    assign coff[3999] = 64'h81665c84ed1f1396;
    assign coff[4000] = 64'h66c0866db3abf1b2;
    assign coff[4001] = 64'h12af33ba815efc65;
    assign coff[4002] = 64'hb3abf1b2993f7993;
    assign coff[4003] = 64'h815efc65ed50cc46;
    assign coff[4004] = 64'h7ea1039bed50cc46;
    assign coff[4005] = 64'h4c540e4e993f7993;
    assign coff[4006] = 64'hed50cc46815efc65;
    assign coff[4007] = 64'h993f7993b3abf1b2;
    assign coff[4008] = 64'h7c23de35e0cda5f5;
    assign coff[4009] = 64'h41b88e849229094f;
    assign coff[4010] = 64'he0cda5f583dc21cb;
    assign coff[4011] = 64'h9229094fbe47717c;
    assign coff[4012] = 64'h6dd6f6b1be47717c;
    assign coff[4013] = 64'h1f325a0b83dc21cb;
    assign coff[4014] = 64'hbe47717c9229094f;
    assign coff[4015] = 64'h83dc21cbe0cda5f5;
    assign coff[4016] = 64'h73ab2ab4c92f28ba;
    assign coff[4017] = 64'h2b078a36877306b4;
    assign coff[4018] = 64'hc92f28ba8c54d54c;
    assign coff[4019] = 64'h877306b4d4f875ca;
    assign coff[4020] = 64'h788cf94cd4f875ca;
    assign coff[4021] = 64'h36d0d7468c54d54c;
    assign coff[4022] = 64'hd4f875ca877306b4;
    assign coff[4023] = 64'h8c54d54cc92f28ba;
    assign coff[4024] = 64'h7fd74964f99f0c68;
    assign coff[4025] = 64'h55e303e6a117a47e;
    assign coff[4026] = 64'hf99f0c688028b69c;
    assign coff[4027] = 64'ha117a47eaa1cfc1a;
    assign coff[4028] = 64'h5ee85b82aa1cfc1a;
    assign coff[4029] = 64'h0660f3988028b69c;
    assign coff[4030] = 64'haa1cfc1aa117a47e;
    assign coff[4031] = 64'h8028b69cf99f0c68;
    assign coff[4032] = 64'h62e20e17aeb8c774;
    assign coff[4033] = 64'h0c72d020809b5541;
    assign coff[4034] = 64'haeb8c7749d1df1e9;
    assign coff[4035] = 64'h809b5541f38d2fe0;
    assign coff[4036] = 64'h7f64aabff38d2fe0;
    assign coff[4037] = 64'h5147388c9d1df1e9;
    assign coff[4038] = 64'hf38d2fe0809b5541;
    assign coff[4039] = 64'h9d1df1e9aeb8c774;
    assign coff[4040] = 64'h7a75b74fdabfe76a;
    assign coff[4041] = 64'h3c408f038f115d72;
    assign coff[4042] = 64'hdabfe76a858a48b1;
    assign coff[4043] = 64'h8f115d72c3bf70fd;
    assign coff[4044] = 64'h70eea28ec3bf70fd;
    assign coff[4045] = 64'h25401896858a48b1;
    assign coff[4046] = 64'hc3bf70fd8f115d72;
    assign coff[4047] = 64'h858a48b1dabfe76a;
    assign coff[4048] = 64'h70d6f0a4c3931c76;
    assign coff[4049] = 64'h250ffeb7857bb152;
    assign coff[4050] = 64'hc3931c768f290f5c;
    assign coff[4051] = 64'h857bb152daf00149;
    assign coff[4052] = 64'h7a844eaedaf00149;
    assign coff[4053] = 64'h3c6ce38a8f290f5c;
    assign coff[4054] = 64'hdaf00149857bb152;
    assign coff[4055] = 64'h8f290f5cc3931c76;
    assign coff[4056] = 64'h7f5fbd77f35b29e0;
    assign coff[4057] = 64'h51205d7b9cfe0e8f;
    assign coff[4058] = 64'hf35b29e080a04289;
    assign coff[4059] = 64'h9cfe0e8faedfa285;
    assign coff[4060] = 64'h6301f171aedfa285;
    assign coff[4061] = 64'h0ca4d62080a04289;
    assign coff[4062] = 64'haedfa2859cfe0e8f;
    assign coff[4063] = 64'h80a04289f35b29e0;
    assign coff[4064] = 64'h6a5fa010b8ce2ecf;
    assign coff[4065] = 64'h18e011678270bbf7;
    assign coff[4066] = 64'hb8ce2ecf95a05ff0;
    assign coff[4067] = 64'h8270bbf7e71fee99;
    assign coff[4068] = 64'h7d8f4409e71fee99;
    assign coff[4069] = 64'h4731d13195a05ff0;
    assign coff[4070] = 64'he71fee998270bbf7;
    assign coff[4071] = 64'h95a05ff0b8ce2ecf;
    assign coff[4072] = 64'h7d85759fe6eea1e4;
    assign coff[4073] = 64'h470805df958472e2;
    assign coff[4074] = 64'he6eea1e4827a8a61;
    assign coff[4075] = 64'h958472e2b8f7fa21;
    assign coff[4076] = 64'h6a7b8d1eb8f7fa21;
    assign coff[4077] = 64'h19115e1c827a8a61;
    assign coff[4078] = 64'hb8f7fa21958472e2;
    assign coff[4079] = 64'h827a8a61e6eea1e4;
    assign coff[4080] = 64'h76380ec8ceed036b;
    assign coff[4081] = 64'h30e48c2289b4b4dd;
    assign coff[4082] = 64'hceed036b89c7f138;
    assign coff[4083] = 64'h89b4b4ddcf1b73de;
    assign coff[4084] = 64'h764b4b23cf1b73de;
    assign coff[4085] = 64'h3112fc9589c7f138;
    assign coff[4086] = 64'hcf1b73de89b4b4dd;
    assign coff[4087] = 64'h89c7f138ceed036b;
    assign coff[4088] = 64'h7ffffd88ffe6de05;
    assign coff[4089] = 64'h5a70b258a56bc2a2;
    assign coff[4090] = 64'hffe6de0580000278;
    assign coff[4091] = 64'ha56bc2a2a58f4da8;
    assign coff[4092] = 64'h5a943d5ea58f4da8;
    assign coff[4093] = 64'h001921fb80000278;
    assign coff[4094] = 64'ha58f4da8a56bc2a2;
    assign coff[4095] = 64'h80000278ffe6de05;
    assign coff[4096] = 64'h5a9d1df1a5983297;
    assign coff[4097] = 64'h0025b2f88000058d;
    assign coff[4098] = 64'ha5983297a562e20f;
    assign coff[4099] = 64'h8000058dffda4d08;
    assign coff[4100] = 64'h7ffffa73ffda4d08;
    assign coff[4101] = 64'h5a67cd69a562e20f;
    assign coff[4102] = 64'hffda4d088000058d;
    assign coff[4103] = 64'ha562e20fa5983297;
    assign coff[4104] = 64'h76501760cf271128;
    assign coff[4105] = 64'h311e978389ccc328;
    assign coff[4106] = 64'hcf27112889afe8a0;
    assign coff[4107] = 64'h89ccc328cee1687d;
    assign coff[4108] = 64'h76333cd8cee1687d;
    assign coff[4109] = 64'h30d8eed889afe8a0;
    assign coff[4110] = 64'hcee1687d89ccc328;
    assign coff[4111] = 64'h89afe8a0cf271128;
    assign coff[4112] = 64'h6a8285d1b9026eac;
    assign coff[4113] = 64'h191db0af827d0102;
    assign coff[4114] = 64'hb9026eac957d7a2f;
    assign coff[4115] = 64'h827d0102e6e24f51;
    assign coff[4116] = 64'h7d82fefee6e24f51;
    assign coff[4117] = 64'h46fd9154957d7a2f;
    assign coff[4118] = 64'he6e24f51827d0102;
    assign coff[4119] = 64'h957d7a2fb9026eac;
    assign coff[4120] = 64'h7d91b49ee72c4260;
    assign coff[4121] = 64'h473c424e95a75dc4;
    assign coff[4122] = 64'he72c4260826e4b62;
    assign coff[4123] = 64'h95a75dc4b8c3bdb2;
    assign coff[4124] = 64'h6a58a23cb8c3bdb2;
    assign coff[4125] = 64'h18d3bda0826e4b62;
    assign coff[4126] = 64'hb8c3bdb295a75dc4;
    assign coff[4127] = 64'h826e4b62e72c4260;
    assign coff[4128] = 64'h6309e7e4aee95b3f;
    assign coff[4129] = 64'h0cb1575280a180ed;
    assign coff[4130] = 64'haee95b3f9cf6181c;
    assign coff[4131] = 64'h80a180edf34ea8ae;
    assign coff[4132] = 64'h7f5e7f13f34ea8ae;
    assign coff[4133] = 64'h5116a4c19cf6181c;
    assign coff[4134] = 64'hf34ea8ae80a180ed;
    assign coff[4135] = 64'h9cf6181caee95b3f;
    assign coff[4136] = 64'h7a87f192dafc08a6;
    assign coff[4137] = 64'h3c77f7378f2efe8f;
    assign coff[4138] = 64'hdafc08a685780e6e;
    assign coff[4139] = 64'h8f2efe8fc38808c9;
    assign coff[4140] = 64'h70d10171c38808c9;
    assign coff[4141] = 64'h2503f75a85780e6e;
    assign coff[4142] = 64'hc38808c98f2efe8f;
    assign coff[4143] = 64'h85780e6edafc08a6;
    assign coff[4144] = 64'h70f48c50c3ca8793;
    assign coff[4145] = 64'h254c1e28858df17c;
    assign coff[4146] = 64'hc3ca87938f0b73b0;
    assign coff[4147] = 64'h858df17cdab3e1d8;
    assign coff[4148] = 64'h7a720e84dab3e1d8;
    assign coff[4149] = 64'h3c35786d8f0b73b0;
    assign coff[4150] = 64'hdab3e1d8858df17c;
    assign coff[4151] = 64'h8f0b73b0c3ca8793;
    assign coff[4152] = 64'h7f65e2fff399b1ad;
    assign coff[4153] = 64'h5150ed5c9d25ed21;
    assign coff[4154] = 64'hf399b1ad809a1d01;
    assign coff[4155] = 64'h9d25ed21aeaf12a4;
    assign coff[4156] = 64'h62da12dfaeaf12a4;
    assign coff[4157] = 64'h0c664e53809a1d01;
    assign coff[4158] = 64'haeaf12a49d25ed21;
    assign coff[4159] = 64'h809a1d01f399b1ad;
    assign coff[4160] = 64'h5ef0c99faa264dce;
    assign coff[4161] = 64'h066d808f8029578b;
    assign coff[4162] = 64'haa264dcea10f3661;
    assign coff[4163] = 64'h8029578bf9927f71;
    assign coff[4164] = 64'h7fd6a875f9927f71;
    assign coff[4165] = 64'h55d9b232a10f3661;
    assign coff[4166] = 64'hf9927f718029578b;
    assign coff[4167] = 64'ha10f3661aa264dce;
    assign coff[4168] = 64'h7891322ad5044bc4;
    assign coff[4169] = 64'h36dc32148c5a3786;
    assign coff[4170] = 64'hd5044bc4876ecdd6;
    assign coff[4171] = 64'h8c5a3786c923cdec;
    assign coff[4172] = 64'h73a5c87ac923cdec;
    assign coff[4173] = 64'h2afbb43c876ecdd6;
    assign coff[4174] = 64'hc923cdec8c5a3786;
    assign coff[4175] = 64'h876ecdd6d5044bc4;
    assign coff[4176] = 64'h6ddd69e9be523a60;
    assign coff[4177] = 64'h1f3e89e083df3273;
    assign coff[4178] = 64'hbe523a6092229617;
    assign coff[4179] = 64'h83df3273e0c17620;
    assign coff[4180] = 64'h7c20cd8de0c17620;
    assign coff[4181] = 64'h41adc5a092229617;
    assign coff[4182] = 64'he0c1762083df3273;
    assign coff[4183] = 64'h92229617be523a60;
    assign coff[4184] = 64'h7ea2d896ed5d3ae5;
    assign coff[4185] = 64'h4c5e24609946f869;
    assign coff[4186] = 64'hed5d3ae5815d276a;
    assign coff[4187] = 64'h9946f869b3a1dba0;
    assign coff[4188] = 64'h66b90797b3a1dba0;
    assign coff[4189] = 64'h12a2c51b815d276a;
    assign coff[4190] = 64'hb3a1dba09946f869;
    assign coff[4191] = 64'h815d276aed5d3ae5;
    assign coff[4192] = 64'h66e5f1beb3de6b17;
    assign coff[4193] = 64'h12ed5a2181683799;
    assign coff[4194] = 64'hb3de6b17991a0e42;
    assign coff[4195] = 64'h81683799ed12a5df;
    assign coff[4196] = 64'h7e97c867ed12a5df;
    assign coff[4197] = 64'h4c2194e9991a0e42;
    assign coff[4198] = 64'hed12a5df81683799;
    assign coff[4199] = 64'h991a0e42b3de6b17;
    assign coff[4200] = 64'h7c331f8ae10a999c;
    assign coff[4201] = 64'h41ee717492495946;
    assign coff[4202] = 64'he10a999c83cce076;
    assign coff[4203] = 64'h92495946be118e8c;
    assign coff[4204] = 64'h6db6a6babe118e8c;
    assign coff[4205] = 64'h1ef5666483cce076;
    assign coff[4206] = 64'hbe118e8c92495946;
    assign coff[4207] = 64'h83cce076e10a999c;
    assign coff[4208] = 64'h73c6051fc967f6ac;
    assign coff[4209] = 64'h2b42b1dd87883477;
    assign coff[4210] = 64'hc967f6ac8c39fae1;
    assign coff[4211] = 64'h87883477d4bd4e23;
    assign coff[4212] = 64'h7877cb89d4bd4e23;
    assign coff[4213] = 64'h369809548c39fae1;
    assign coff[4214] = 64'hd4bd4e2387883477;
    assign coff[4215] = 64'h8c39fae1c967f6ac;
    assign coff[4216] = 64'h7fda5b8ff9ddce22;
    assign coff[4217] = 64'h56118ffea141d8c5;
    assign coff[4218] = 64'hf9ddce228025a471;
    assign coff[4219] = 64'ha141d8c5a9ee7002;
    assign coff[4220] = 64'h5ebe273ba9ee7002;
    assign coff[4221] = 64'h062231de8025a471;
    assign coff[4222] = 64'ha9ee7002a141d8c5;
    assign coff[4223] = 64'h8025a471f9ddce22;
    assign coff[4224] = 64'h5cce1b97a7d8742f;
    assign coff[4225] = 64'h0349daac800ad0e3;
    assign coff[4226] = 64'ha7d8742fa331e469;
    assign coff[4227] = 64'h800ad0e3fcb62554;
    assign coff[4228] = 64'h7ff52f1dfcb62554;
    assign coff[4229] = 64'h58278bd1a331e469;
    assign coff[4230] = 64'hfcb62554800ad0e3;
    assign coff[4231] = 64'ha331e469a7d8742f;
    assign coff[4232] = 64'h7779db03d21223e7;
    assign coff[4233] = 64'h3401674a8b0a78c7;
    assign coff[4234] = 64'hd21223e7888624fd;
    assign coff[4235] = 64'h8b0a78c7cbfe98b6;
    assign coff[4236] = 64'h74f58739cbfe98b6;
    assign coff[4237] = 64'h2deddc19888624fd;
    assign coff[4238] = 64'hcbfe98b68b0a78c7;
    assign coff[4239] = 64'h888624fdd21223e7;
    assign coff[4240] = 64'h6c384fefbba50f50;
    assign coff[4241] = 64'h1c3049ac83247943;
    assign coff[4242] = 64'hbba50f5093c7b011;
    assign coff[4243] = 64'h83247943e3cfb654;
    assign coff[4244] = 64'h7cdb86bde3cfb654;
    assign coff[4245] = 64'h445af0b093c7b011;
    assign coff[4246] = 64'he3cfb65483247943;
    assign coff[4247] = 64'h93c7b011bba50f50;
    assign coff[4248] = 64'h7e240064ea431191;
    assign coff[4249] = 64'h49d2e47e976f1b24;
    assign coff[4250] = 64'hea43119181dbff9c;
    assign coff[4251] = 64'h976f1b24b62d1b82;
    assign coff[4252] = 64'h6890e4dcb62d1b82;
    assign coff[4253] = 64'h15bcee6f81dbff9c;
    assign coff[4254] = 64'hb62d1b82976f1b24;
    assign coff[4255] = 64'h81dbff9cea431191;
    assign coff[4256] = 64'h64ffb65bb15dd315;
    assign coff[4257] = 64'h0fd090e180fb1121;
    assign coff[4258] = 64'hb15dd3159b0049a5;
    assign coff[4259] = 64'h80fb1121f02f6f1f;
    assign coff[4260] = 64'h7f04eedff02f6f1f;
    assign coff[4261] = 64'h4ea22ceb9b0049a5;
    assign coff[4262] = 64'hf02f6f1f80fb1121;
    assign coff[4263] = 64'h9b0049a5b15dd315;
    assign coff[4264] = 64'h7b670c4dde00b216;
    assign coff[4265] = 64'h3f38142a90b39715;
    assign coff[4266] = 64'hde00b2168498f3b3;
    assign coff[4267] = 64'h90b39715c0c7ebd6;
    assign coff[4268] = 64'h6f4c68ebc0c7ebd6;
    assign coff[4269] = 64'h21ff4dea8498f3b3;
    assign coff[4270] = 64'hc0c7ebd690b39715;
    assign coff[4271] = 64'h8498f3b3de00b216;
    assign coff[4272] = 64'h72661abfc694d1c8;
    assign coff[4273] = 64'h284a83498681b4ea;
    assign coff[4274] = 64'hc694d1c88d99e541;
    assign coff[4275] = 64'h8681b4ead7b57cb7;
    assign coff[4276] = 64'h797e4b16d7b57cb7;
    assign coff[4277] = 64'h396b2e388d99e541;
    assign coff[4278] = 64'hd7b57cb78681b4ea;
    assign coff[4279] = 64'h8d99e541c694d1c8;
    assign coff[4280] = 64'h7fa9f723f6bb08f1;
    assign coff[4281] = 64'h53b7b31c9f2c6bc5;
    assign coff[4282] = 64'hf6bb08f1805608dd;
    assign coff[4283] = 64'h9f2c6bc5ac484ce4;
    assign coff[4284] = 64'h60d3943bac484ce4;
    assign coff[4285] = 64'h0944f70f805608dd;
    assign coff[4286] = 64'hac484ce49f2c6bc5;
    assign coff[4287] = 64'h805608ddf6bb08f1;
    assign coff[4288] = 64'h6104d3bcac81647e;
    assign coff[4289] = 64'h099028b3805b94ce;
    assign coff[4290] = 64'hac81647e9efb2c44;
    assign coff[4291] = 64'h805b94cef66fd74d;
    assign coff[4292] = 64'h7fa46b32f66fd74d;
    assign coff[4293] = 64'h537e9b829efb2c44;
    assign coff[4294] = 64'hf66fd74d805b94ce;
    assign coff[4295] = 64'h9efb2c44ac81647e;
    assign coff[4296] = 64'h7995f1c1d7fd1474;
    assign coff[4297] = 64'h39ae872f8dbbcba0;
    assign coff[4298] = 64'hd7fd1474866a0e3f;
    assign coff[4299] = 64'h8dbbcba0c65178d1;
    assign coff[4300] = 64'h72443460c65178d1;
    assign coff[4301] = 64'h2802eb8c866a0e3f;
    assign coff[4302] = 64'hc65178d18dbbcba0;
    assign coff[4303] = 64'h866a0e3fd7fd1474;
    assign coff[4304] = 64'h6f7192cfc1098634;
    assign coff[4305] = 64'h2247f8aa84ad0fc6;
    assign coff[4306] = 64'hc1098634908e6d31;
    assign coff[4307] = 64'h84ad0fc6ddb80756;
    assign coff[4308] = 64'h7b52f03addb80756;
    assign coff[4309] = 64'h3ef679cc908e6d31;
    assign coff[4310] = 64'hddb8075684ad0fc6;
    assign coff[4311] = 64'h908e6d31c1098634;
    assign coff[4312] = 64'h7f0e29a3f07a43e7;
    assign coff[4313] = 64'h4edd9d899b2eaccf;
    assign coff[4314] = 64'hf07a43e780f1d65d;
    assign coff[4315] = 64'h9b2eaccfb1226277;
    assign coff[4316] = 64'h64d15331b1226277;
    assign coff[4317] = 64'h0f85bc1980f1d65d;
    assign coff[4318] = 64'hb12262779b2eaccf;
    assign coff[4319] = 64'h80f1d65df07a43e7;
    assign coff[4320] = 64'h68bc4f13b66ac07c;
    assign coff[4321] = 64'h1607383481e8e381;
    assign coff[4322] = 64'hb66ac07c9743b0ed;
    assign coff[4323] = 64'h81e8e381e9f8c7cc;
    assign coff[4324] = 64'h7e171c7fe9f8c7cc;
    assign coff[4325] = 64'h49953f849743b0ed;
    assign coff[4326] = 64'he9f8c7cc81e8e381;
    assign coff[4327] = 64'h9743b0edb66ac07c;
    assign coff[4328] = 64'h7cec0bd1e4194746;
    assign coff[4329] = 64'h449aa40093f0068f;
    assign coff[4330] = 64'he41947468313f42f;
    assign coff[4331] = 64'h93f0068fbb655c00;
    assign coff[4332] = 64'h6c0ff971bb655c00;
    assign coff[4333] = 64'h1be6b8ba8313f42f;
    assign coff[4334] = 64'hbb655c0093f0068f;
    assign coff[4335] = 64'h8313f42fe4194746;
    assign coff[4336] = 64'h7514152bcc4386bc;
    assign coff[4337] = 64'h2e3434ac88a147a9;
    assign coff[4338] = 64'hcc4386bc8aebead5;
    assign coff[4339] = 64'h88a147a9d1cbcb54;
    assign coff[4340] = 64'h775eb857d1cbcb54;
    assign coff[4341] = 64'h33bc79448aebead5;
    assign coff[4342] = 64'hd1cbcb5488a147a9;
    assign coff[4343] = 64'h8aebead5cc4386bc;
    assign coff[4344] = 64'h7ff708cefd018574;
    assign coff[4345] = 64'h585e2730a365e1e2;
    assign coff[4346] = 64'hfd0185748008f732;
    assign coff[4347] = 64'ha365e1e2a7a1d8d0;
    assign coff[4348] = 64'h5c9a1e1ea7a1d8d0;
    assign coff[4349] = 64'h02fe7a8c8008f732;
    assign coff[4350] = 64'ha7a1d8d0a365e1e2;
    assign coff[4351] = 64'h8008f732fd018574;
    assign coff[4352] = 64'h5bb7615da6b69ac8;
    assign coff[4353] = 64'h01b7cf4d8002f3a1;
    assign coff[4354] = 64'ha6b69ac8a4489ea3;
    assign coff[4355] = 64'h8002f3a1fe4830b3;
    assign coff[4356] = 64'h7ffd0c5ffe4830b3;
    assign coff[4357] = 64'h59496538a4489ea3;
    assign coff[4358] = 64'hfe4830b38002f3a1;
    assign coff[4359] = 64'ha4489ea3a6b69ac8;
    assign coff[4360] = 64'h76e743f4d09bb0aa;
    assign coff[4361] = 64'h3290f8ef8a6959b3;
    assign coff[4362] = 64'hd09bb0aa8918bc0c;
    assign coff[4363] = 64'h8a6959b3cd6f0711;
    assign coff[4364] = 64'h7596a64dcd6f0711;
    assign coff[4365] = 64'h2f644f568918bc0c;
    assign coff[4366] = 64'hcd6f07118a6959b3;
    assign coff[4367] = 64'h8918bc0cd09bb0aa;
    assign coff[4368] = 64'h6b5f7cbcba526726;
    assign coff[4369] = 64'h1aa780b682ce5356;
    assign coff[4370] = 64'hba52672694a08344;
    assign coff[4371] = 64'h82ce5356e5587f4a;
    assign coff[4372] = 64'h7d31acaae5587f4a;
    assign coff[4373] = 64'h45ad98da94a08344;
    assign coff[4374] = 64'he5587f4a82ce5356;
    assign coff[4375] = 64'h94a08344ba526726;
    assign coff[4376] = 64'h7ddd479de8b73712;
    assign coff[4377] = 64'h4888f95796893404;
    assign coff[4378] = 64'he8b737128222b863;
    assign coff[4379] = 64'h96893404b77706a9;
    assign coff[4380] = 64'h6976cbfcb77706a9;
    assign coff[4381] = 64'h1748c8ee8222b863;
    assign coff[4382] = 64'hb77706a996893404;
    assign coff[4383] = 64'h8222b863e8b73712;
    assign coff[4384] = 64'h6406bcbab0220d0a;
    assign coff[4385] = 64'h0e413a7280cbd54f;
    assign coff[4386] = 64'hb0220d0a9bf94346;
    assign coff[4387] = 64'h80cbd54ff1bec58e;
    assign coff[4388] = 64'h7f342ab1f1bec58e;
    assign coff[4389] = 64'h4fddf2f69bf94346;
    assign coff[4390] = 64'hf1bec58e80cbd54f;
    assign coff[4391] = 64'h9bf94346b0220d0a;
    assign coff[4392] = 64'h7af9ddcbdc7dae23;
    assign coff[4393] = 64'h3dd936e68fef21ce;
    assign coff[4394] = 64'hdc7dae2385062235;
    assign coff[4395] = 64'h8fef21cec226c91a;
    assign coff[4396] = 64'h7010de32c226c91a;
    assign coff[4397] = 64'h238251dd85062235;
    assign coff[4398] = 64'hc226c91a8fef21ce;
    assign coff[4399] = 64'h85062235dc7dae23;
    assign coff[4400] = 64'h71af848ac52e8a6d;
    assign coff[4401] = 64'h26cc102d86057944;
    assign coff[4402] = 64'hc52e8a6d8e507b76;
    assign coff[4403] = 64'h86057944d933efd3;
    assign coff[4404] = 64'h79fa86bcd933efd3;
    assign coff[4405] = 64'h3ad175938e507b76;
    assign coff[4406] = 64'hd933efd386057944;
    assign coff[4407] = 64'h8e507b76c52e8a6d;
    assign coff[4408] = 64'h7f8a6272f52a27d7;
    assign coff[4409] = 64'h5285e7779e27499a;
    assign coff[4410] = 64'hf52a27d780759d8e;
    assign coff[4411] = 64'h9e27499aad7a1889;
    assign coff[4412] = 64'h61d8b666ad7a1889;
    assign coff[4413] = 64'h0ad5d82980759d8e;
    assign coff[4414] = 64'had7a18899e27499a;
    assign coff[4415] = 64'h80759d8ef52a27d7;
    assign coff[4416] = 64'h5ffca859ab523748;
    assign coff[4417] = 64'h07fefc16803fffc2;
    assign coff[4418] = 64'hab523748a00357a7;
    assign coff[4419] = 64'h803fffc2f80103ea;
    assign coff[4420] = 64'h7fc0003ef80103ea;
    assign coff[4421] = 64'h54adc8b8a00357a7;
    assign coff[4422] = 64'hf80103ea803fffc2;
    assign coff[4423] = 64'ha00357a7ab523748;
    assign coff[4424] = 64'h7915e77cd67fe351;
    assign coff[4425] = 64'h384672558d08ca40;
    assign coff[4426] = 64'hd67fe35186ea1884;
    assign coff[4427] = 64'h8d08ca40c7b98dab;
    assign coff[4428] = 64'h72f735c0c7b98dab;
    assign coff[4429] = 64'h29801caf86ea1884;
    assign coff[4430] = 64'hc7b98dab8d08ca40;
    assign coff[4431] = 64'h86ea1884d67fe351;
    assign coff[4432] = 64'h6ea9a073bfaca2dc;
    assign coff[4433] = 64'h20c3e2f58443be82;
    assign coff[4434] = 64'hbfaca2dc91565f8d;
    assign coff[4435] = 64'h8443be82df3c1d0b;
    assign coff[4436] = 64'h7bbc417edf3c1d0b;
    assign coff[4437] = 64'h40535d2491565f8d;
    assign coff[4438] = 64'hdf3c1d0b8443be82;
    assign coff[4439] = 64'h91565f8dbfaca2dc;
    assign coff[4440] = 64'h7edaf31ceeeb6b1c;
    assign coff[4441] = 64'h4d9f60019a38dc5d;
    assign coff[4442] = 64'heeeb6b1c81250ce4;
    assign coff[4443] = 64'h9a38dc5db2609fff;
    assign coff[4444] = 64'h65c723a3b2609fff;
    assign coff[4445] = 64'h111494e481250ce4;
    assign coff[4446] = 64'hb2609fff9a38dc5d;
    assign coff[4447] = 64'h81250ce4eeeb6b1c;
    assign coff[4448] = 64'h67d320c1b523245b;
    assign coff[4449] = 64'h147aae3a81a61e0b;
    assign coff[4450] = 64'hb523245b982cdf3f;
    assign coff[4451] = 64'h81a61e0beb8551c6;
    assign coff[4452] = 64'h7e59e1f5eb8551c6;
    assign coff[4453] = 64'h4adcdba5982cdf3f;
    assign coff[4454] = 64'heb8551c681a61e0b;
    assign coff[4455] = 64'h982cdf3fb523245b;
    assign coff[4456] = 64'h7c91fc66e2915f34;
    assign coff[4457] = 64'h4345d6b3931a968b;
    assign coff[4458] = 64'he2915f34836e039a;
    assign coff[4459] = 64'h931a968bbcba294d;
    assign coff[4460] = 64'h6ce56975bcba294d;
    assign coff[4461] = 64'h1d6ea0cc836e039a;
    assign coff[4462] = 64'hbcba294d931a968b;
    assign coff[4463] = 64'h836e039ae2915f34;
    assign coff[4464] = 64'h746f4bb8cad4b853;
    assign coff[4465] = 64'h2cbc500688126e40;
    assign coff[4466] = 64'hcad4b8538b90b448;
    assign coff[4467] = 64'h88126e40d343affa;
    assign coff[4468] = 64'h77ed91c0d343affa;
    assign coff[4469] = 64'h352b47ad8b90b448;
    assign coff[4470] = 64'hd343affa88126e40;
    assign coff[4471] = 64'h8b90b448cad4b853;
    assign coff[4472] = 64'h7feb296dfb6f9345;
    assign coff[4473] = 64'h57398a05a2520f0b;
    assign coff[4474] = 64'hfb6f93458014d693;
    assign coff[4475] = 64'ha2520f0ba8c675fb;
    assign coff[4476] = 64'h5dadf0f5a8c675fb;
    assign coff[4477] = 64'h04906cbb8014d693;
    assign coff[4478] = 64'ha8c675fba2520f0b;
    assign coff[4479] = 64'h8014d693fb6f9345;
    assign coff[4480] = 64'h5de141e1a8fdb3a1;
    assign coff[4481] = 64'h04dbc59780179d06;
    assign coff[4482] = 64'ha8fdb3a1a21ebe1f;
    assign coff[4483] = 64'h80179d06fb243a69;
    assign coff[4484] = 64'h7fe862fafb243a69;
    assign coff[4485] = 64'h57024c5fa21ebe1f;
    assign coff[4486] = 64'hfb243a6980179d06;
    assign coff[4487] = 64'ha21ebe1fa8fdb3a1;
    assign coff[4488] = 64'h7807d6e9d38a5c70;
    assign coff[4489] = 64'h356fd4618bb01a2e;
    assign coff[4490] = 64'hd38a5c7087f82917;
    assign coff[4491] = 64'h8bb01a2eca902b9f;
    assign coff[4492] = 64'h744fe5d2ca902b9f;
    assign coff[4493] = 64'h2c75a39087f82917;
    assign coff[4494] = 64'hca902b9f8bb01a2e;
    assign coff[4495] = 64'h87f82917d38a5c70;
    assign coff[4496] = 64'h6d0cf70fbcfa5a1b;
    assign coff[4497] = 64'h1db7fc6d837f6f78;
    assign coff[4498] = 64'hbcfa5a1b92f308f1;
    assign coff[4499] = 64'h837f6f78e2480393;
    assign coff[4500] = 64'h7c809088e2480393;
    assign coff[4501] = 64'h4305a5e592f308f1;
    assign coff[4502] = 64'he2480393837f6f78;
    assign coff[4503] = 64'h92f308f1bcfa5a1b;
    assign coff[4504] = 64'h7e65dc3bebcfc29b;
    assign coff[4505] = 64'h4b19f70a98590a48;
    assign coff[4506] = 64'hebcfc29b819a23c5;
    assign coff[4507] = 64'h98590a48b4e608f6;
    assign coff[4508] = 64'h67a6f5b8b4e608f6;
    assign coff[4509] = 64'h14303d65819a23c5;
    assign coff[4510] = 64'hb4e608f698590a48;
    assign coff[4511] = 64'h819a23c5ebcfc29b;
    assign coff[4512] = 64'h65f4cb2db29ca132;
    assign coff[4513] = 64'h115f4b3c812f3290;
    assign coff[4514] = 64'hb29ca1329a0b34d3;
    assign coff[4515] = 64'h812f3290eea0b4c4;
    assign coff[4516] = 64'h7ed0cd70eea0b4c4;
    assign coff[4517] = 64'h4d635ece9a0b34d3;
    assign coff[4518] = 64'heea0b4c4812f3290;
    assign coff[4519] = 64'h9a0b34d3b29ca132;
    assign coff[4520] = 64'h7bcf78e5df850591;
    assign coff[4521] = 64'h4094817f917c56d1;
    assign coff[4522] = 64'hdf8505918430871b;
    assign coff[4523] = 64'h917c56d1bf6b7e81;
    assign coff[4524] = 64'h6e83a92fbf6b7e81;
    assign coff[4525] = 64'h207afa6f8430871b;
    assign coff[4526] = 64'hbf6b7e81917c56d1;
    assign coff[4527] = 64'h8430871bdf850591;
    assign coff[4528] = 64'h731847e5c7fd4fd4;
    assign coff[4529] = 64'h29c768be87029fa3;
    assign coff[4530] = 64'hc7fd4fd48ce7b81b;
    assign coff[4531] = 64'h87029fa3d6389742;
    assign coff[4532] = 64'h78fd605dd6389742;
    assign coff[4533] = 64'h3802b02c8ce7b81b;
    assign coff[4534] = 64'hd638974287029fa3;
    assign coff[4535] = 64'h8ce7b81bc7fd4fd4;
    assign coff[4536] = 64'h7fc49fdaf84c4588;
    assign coff[4537] = 64'h54e64482a0354990;
    assign coff[4538] = 64'hf84c4588803b6026;
    assign coff[4539] = 64'ha0354990ab19bb7e;
    assign coff[4540] = 64'h5fcab670ab19bb7e;
    assign coff[4541] = 64'h07b3ba78803b6026;
    assign coff[4542] = 64'hab19bb7ea0354990;
    assign coff[4543] = 64'h803b6026f84c4588;
    assign coff[4544] = 64'h62094199adb3c9c0;
    assign coff[4545] = 64'h0b20f6ee807c159c;
    assign coff[4546] = 64'hadb3c9c09df6be67;
    assign coff[4547] = 64'h807c159cf4df0912;
    assign coff[4548] = 64'h7f83ea64f4df0912;
    assign coff[4549] = 64'h524c36409df6be67;
    assign coff[4550] = 64'hf4df0912807c159c;
    assign coff[4551] = 64'h9df6be67adb3c9c0;
    assign coff[4552] = 64'h7a114c09d97bd07c;
    assign coff[4553] = 64'h3b1462be8e7334c1;
    assign coff[4554] = 64'hd97bd07c85eeb3f7;
    assign coff[4555] = 64'h8e7334c1c4eb9d42;
    assign coff[4556] = 64'h718ccb3fc4eb9d42;
    assign coff[4557] = 64'h26842f8485eeb3f7;
    assign coff[4558] = 64'hc4eb9d428e7334c1;
    assign coff[4559] = 64'h85eeb3f7d97bd07c;
    assign coff[4560] = 64'h70353947c268d6f5;
    assign coff[4561] = 64'h23cabc09851b222e;
    assign coff[4562] = 64'hc268d6f58fcac6b9;
    assign coff[4563] = 64'h851b222edc3543f7;
    assign coff[4564] = 64'h7ae4ddd2dc3543f7;
    assign coff[4565] = 64'h3d97290b8fcac6b9;
    assign coff[4566] = 64'hdc3543f7851b222e;
    assign coff[4567] = 64'h8fcac6b9c268d6f5;
    assign coff[4568] = 64'h7f3c7a31f209b5e4;
    assign coff[4569] = 64'h5018d0b49c286046;
    assign coff[4570] = 64'hf209b5e480c385cf;
    assign coff[4571] = 64'h9c286046afe72f4c;
    assign coff[4572] = 64'h63d79fbaafe72f4c;
    assign coff[4573] = 64'h0df64a1c80c385cf;
    assign coff[4574] = 64'hafe72f4c9c286046;
    assign coff[4575] = 64'h80c385cff209b5e4;
    assign coff[4576] = 64'h69a173b5b7b532d6;
    assign coff[4577] = 64'h1792e8c68230856a;
    assign coff[4578] = 64'hb7b532d6965e8c4b;
    assign coff[4579] = 64'h8230856ae86d173a;
    assign coff[4580] = 64'h7dcf7a96e86d173a;
    assign coff[4581] = 64'h484acd2a965e8c4b;
    assign coff[4582] = 64'he86d173a8230856a;
    assign coff[4583] = 64'h965e8c4bb7b532d6;
    assign coff[4584] = 64'h7d414a51e5a242b7;
    assign coff[4585] = 64'h45eccc3794c9a119;
    assign coff[4586] = 64'he5a242b782beb5af;
    assign coff[4587] = 64'h94c9a119ba1333c9;
    assign coff[4588] = 64'h6b365ee7ba1333c9;
    assign coff[4589] = 64'h1a5dbd4982beb5af;
    assign coff[4590] = 64'hba1333c994c9a119;
    assign coff[4591] = 64'h82beb5afe5a242b7;
    assign coff[4592] = 64'h75b45b1dcdb453c0;
    assign coff[4593] = 64'h2faa514f8934bb31;
    assign coff[4594] = 64'hcdb453c08a4ba4e3;
    assign coff[4595] = 64'h8934bb31d055aeb1;
    assign coff[4596] = 64'h76cb44cfd055aeb1;
    assign coff[4597] = 64'h324bac408a4ba4e3;
    assign coff[4598] = 64'hd055aeb18934bb31;
    assign coff[4599] = 64'h8a4ba4e3cdb453c0;
    assign coff[4600] = 64'h7ffdf93cfe939530;
    assign coff[4601] = 64'h597f5c36a47d46a8;
    assign coff[4602] = 64'hfe939530800206c4;
    assign coff[4603] = 64'ha47d46a8a680a3ca;
    assign coff[4604] = 64'h5b82b958a680a3ca;
    assign coff[4605] = 64'h016c6ad0800206c4;
    assign coff[4606] = 64'ha680a3caa47d46a8;
    assign coff[4607] = 64'h800206c4fe939530;
    assign coff[4608] = 64'h5b2ab020a626f7d7;
    assign coff[4609] = 64'h00eec2498000deaf;
    assign coff[4610] = 64'ha626f7d7a4d54fe0;
    assign coff[4611] = 64'h8000deafff113db7;
    assign coff[4612] = 64'h7fff2151ff113db7;
    assign coff[4613] = 64'h59d90829a4d54fe0;
    assign coff[4614] = 64'hff113db78000deaf;
    assign coff[4615] = 64'ha4d54fe0a626f7d7;
    assign coff[4616] = 64'h769c3ffecfe1258b;
    assign coff[4617] = 64'h31d805b78a1a7cfb;
    assign coff[4618] = 64'hcfe1258b8963c002;
    assign coff[4619] = 64'h8a1a7cfbce27fa49;
    assign coff[4620] = 64'h75e58305ce27fa49;
    assign coff[4621] = 64'h301eda758963c002;
    assign coff[4622] = 64'hce27fa498a1a7cfb;
    assign coff[4623] = 64'h8963c002cfe1258b;
    assign coff[4624] = 64'h6af18536b9aa1423;
    assign coff[4625] = 64'h19e2b8a282a50f85;
    assign coff[4626] = 64'hb9aa1423950e7aca;
    assign coff[4627] = 64'h82a50f85e61d475e;
    assign coff[4628] = 64'h7d5af07be61d475e;
    assign coff[4629] = 64'h4655ebdd950e7aca;
    assign coff[4630] = 64'he61d475e82a50f85;
    assign coff[4631] = 64'h950e7acab9aa1423;
    assign coff[4632] = 64'h7db81936e7f19f0c;
    assign coff[4633] = 64'h47e2f6829617c63c;
    assign coff[4634] = 64'he7f19f0c8247e6ca;
    assign coff[4635] = 64'h9617c63cb81d097e;
    assign coff[4636] = 64'h69e839c4b81d097e;
    assign coff[4637] = 64'h180e60f48247e6ca;
    assign coff[4638] = 64'hb81d097e9617c63c;
    assign coff[4639] = 64'h8247e6cae7f19f0c;
    assign coff[4640] = 64'h6388cd1baf8550db;
    assign coff[4641] = 64'h0d79598280b60e15;
    assign coff[4642] = 64'haf8550db9c7732e5;
    assign coff[4643] = 64'h80b60e15f286a67e;
    assign coff[4644] = 64'h7f49f1ebf286a67e;
    assign coff[4645] = 64'h507aaf259c7732e5;
    assign coff[4646] = 64'hf286a67e80b60e15;
    assign coff[4647] = 64'h9c7732e5af8550db;
    assign coff[4648] = 64'h7ac17f20dbbcaea8;
    assign coff[4649] = 64'h3d28e2828f8e8576;
    assign coff[4650] = 64'hdbbcaea8853e80e0;
    assign coff[4651] = 64'h8f8e8576c2d71d7e;
    assign coff[4652] = 64'h70717a8ac2d71d7e;
    assign coff[4653] = 64'h24435158853e80e0;
    assign coff[4654] = 64'hc2d71d7e8f8e8576;
    assign coff[4655] = 64'h853e80e0dbbcaea8;
    assign coff[4656] = 64'h7152943bc47c3f94;
    assign coff[4657] = 64'h260c461b85c91e9a;
    assign coff[4658] = 64'hc47c3f948ead6bc5;
    assign coff[4659] = 64'h85c91e9ad9f3b9e5;
    assign coff[4660] = 64'h7a36e166d9f3b9e5;
    assign coff[4661] = 64'h3b83c06c8ead6bc5;
    assign coff[4662] = 64'hd9f3b9e585c91e9a;
    assign coff[4663] = 64'h8ead6bc5c47c3f94;
    assign coff[4664] = 64'h7f78bffbf461de6d;
    assign coff[4665] = 64'h51ebcf7a9da62208;
    assign coff[4666] = 64'hf461de6d80874005;
    assign coff[4667] = 64'h9da62208ae143086;
    assign coff[4668] = 64'h6259ddf8ae143086;
    assign coff[4669] = 64'h0b9e219380874005;
    assign coff[4670] = 64'hae1430869da62208;
    assign coff[4671] = 64'h80874005f461de6d;
    assign coff[4672] = 64'h5f772ec2aabbd959;
    assign coff[4673] = 64'h0736473880340dfd;
    assign coff[4674] = 64'haabbd959a088d13e;
    assign coff[4675] = 64'h80340dfdf8c9b8c8;
    assign coff[4676] = 64'h7fcbf203f8c9b8c8;
    assign coff[4677] = 64'h554426a7a088d13e;
    assign coff[4678] = 64'hf8c9b8c880340dfd;
    assign coff[4679] = 64'ha088d13eaabbd959;
    assign coff[4680] = 64'h78d421e4d5c1e36d;
    assign coff[4681] = 64'h379196c38cb0f2a1;
    assign coff[4682] = 64'hd5c1e36d872bde1c;
    assign coff[4683] = 64'h8cb0f2a1c86e693d;
    assign coff[4684] = 64'h734f0d5fc86e693d;
    assign coff[4685] = 64'h2a3e1c93872bde1c;
    assign coff[4686] = 64'hc86e693d8cb0f2a1;
    assign coff[4687] = 64'h872bde1cd5c1e36d;
    assign coff[4688] = 64'h6e440d37beff1e6c;
    assign coff[4689] = 64'h20015de78410df95;
    assign coff[4690] = 64'hbeff1e6c91bbf2c9;
    assign coff[4691] = 64'h8410df95dffea219;
    assign coff[4692] = 64'h7bef206bdffea219;
    assign coff[4693] = 64'h4100e19491bbf2c9;
    assign coff[4694] = 64'hdffea2198410df95;
    assign coff[4695] = 64'h91bbf2c9beff1e6c;
    assign coff[4696] = 64'h7ebf8237ee243cf9;
    assign coff[4697] = 64'h4cff212e99bf6c3d;
    assign coff[4698] = 64'hee243cf981407dc9;
    assign coff[4699] = 64'h99bf6c3db300ded2;
    assign coff[4700] = 64'h664093c3b300ded2;
    assign coff[4701] = 64'h11dbc30781407dc9;
    assign coff[4702] = 64'hb300ded299bf6c3d;
    assign coff[4703] = 64'h81407dc9ee243cf9;
    assign coff[4704] = 64'h675d08c4b4806a95;
    assign coff[4705] = 64'h13b41c7d81868eca;
    assign coff[4706] = 64'hb4806a9598a2f73c;
    assign coff[4707] = 64'h81868ecaec4be383;
    assign coff[4708] = 64'h7e797136ec4be383;
    assign coff[4709] = 64'h4b7f956b98a2f73c;
    assign coff[4710] = 64'hec4be38381868eca;
    assign coff[4711] = 64'h98a2f73cb4806a95;
    assign coff[4712] = 64'h7c63276de1cdd727;
    assign coff[4713] = 64'h429a763f92b1710e;
    assign coff[4714] = 64'he1cdd727839cd893;
    assign coff[4715] = 64'h92b1710ebd6589c1;
    assign coff[4716] = 64'h6d4e8ef2bd6589c1;
    assign coff[4717] = 64'h1e3228d9839cd893;
    assign coff[4718] = 64'hbd6589c192b1710e;
    assign coff[4719] = 64'h839cd893e1cdd727;
    assign coff[4720] = 64'h741b37a9ca1e1506;
    assign coff[4721] = 64'h2bffb73a87ccbd11;
    assign coff[4722] = 64'hca1e15068be4c857;
    assign coff[4723] = 64'h87ccbd11d40048c6;
    assign coff[4724] = 64'h783342efd40048c6;
    assign coff[4725] = 64'h35e1eafa8be4c857;
    assign coff[4726] = 64'hd40048c687ccbd11;
    assign coff[4727] = 64'h8be4c857ca1e1506;
    assign coff[4728] = 64'h7fe36045faa6aa1a;
    assign coff[4729] = 64'h56a5f7e7a1c97fad;
    assign coff[4730] = 64'hfaa6aa1a801c9fbb;
    assign coff[4731] = 64'ha1c97fada95a0819;
    assign coff[4732] = 64'h5e368053a95a0819;
    assign coff[4733] = 64'h055955e6801c9fbb;
    assign coff[4734] = 64'ha95a0819a1c97fad;
    assign coff[4735] = 64'h801c9fbbfaa6aa1a;
    assign coff[4736] = 64'h5d5821e4a86aa7db;
    assign coff[4737] = 64'h0412d5288010991f;
    assign coff[4738] = 64'ha86aa7dba2a7de1c;
    assign coff[4739] = 64'h8010991ffbed2ad8;
    assign coff[4740] = 64'h7fef66e1fbed2ad8;
    assign coff[4741] = 64'h57955825a2a7de1c;
    assign coff[4742] = 64'hfbed2ad88010991f;
    assign coff[4743] = 64'ha2a7de1ca86aa7db;
    assign coff[4744] = 64'h77c16cb4d2ce0869;
    assign coff[4745] = 64'h34b8dee18b5cb995;
    assign coff[4746] = 64'hd2ce0869883e934c;
    assign coff[4747] = 64'h8b5cb995cb47211f;
    assign coff[4748] = 64'h74a3466bcb47211f;
    assign coff[4749] = 64'h2d31f797883e934c;
    assign coff[4750] = 64'hcb47211f8b5cb995;
    assign coff[4751] = 64'h883e934cd2ce0869;
    assign coff[4752] = 64'h6ca32985bc4f6134;
    assign coff[4753] = 64'h1cf446c583515a8c;
    assign coff[4754] = 64'hbc4f6134935cd67b;
    assign coff[4755] = 64'h83515a8ce30bb93b;
    assign coff[4756] = 64'h7caea574e30bb93b;
    assign coff[4757] = 64'h43b09ecc935cd67b;
    assign coff[4758] = 64'he30bb93b83515a8c;
    assign coff[4759] = 64'h935cd67bbc4f6134;
    assign coff[4760] = 64'h7e458a17eb095039;
    assign coff[4761] = 64'h4a76c9a297e39245;
    assign coff[4762] = 64'heb09503981ba75e9;
    assign coff[4763] = 64'h97e39245b589365e;
    assign coff[4764] = 64'h681c6dbbb589365e;
    assign coff[4765] = 64'h14f6afc781ba75e9;
    assign coff[4766] = 64'hb589365e97e39245;
    assign coff[4767] = 64'h81ba75e9eb095039;
    assign coff[4768] = 64'h657abdf6b1fcd9e5;
    assign coff[4769] = 64'h1098028781148544;
    assign coff[4770] = 64'hb1fcd9e59a85420a;
    assign coff[4771] = 64'h81148544ef67fd79;
    assign coff[4772] = 64'h7eeb7abcef67fd79;
    assign coff[4773] = 64'h4e03261b9a85420a;
    assign coff[4774] = 64'hef67fd7981148544;
    assign coff[4775] = 64'h9a85420ab1fcd9e5;
    assign coff[4776] = 64'h7b9bdb18dec2b2d1;
    assign coff[4777] = 64'h3fe699aa91176e1f;
    assign coff[4778] = 64'hdec2b2d1846424e8;
    assign coff[4779] = 64'h91176e1fc0196656;
    assign coff[4780] = 64'h6ee891e1c0196656;
    assign coff[4781] = 64'h213d4d2f846424e8;
    assign coff[4782] = 64'hc019665691176e1f;
    assign coff[4783] = 64'h846424e8dec2b2d1;
    assign coff[4784] = 64'h72bfbee3c748cad6;
    assign coff[4785] = 64'h290928a386c194b2;
    assign coff[4786] = 64'hc748cad68d40411d;
    assign coff[4787] = 64'h86c194b2d6f6d75d;
    assign coff[4788] = 64'h793e6b4ed6f6d75d;
    assign coff[4789] = 64'h38b7352a8d40411d;
    assign coff[4790] = 64'hd6f6d75d86c194b2;
    assign coff[4791] = 64'h8d40411dc748cad6;
    assign coff[4792] = 64'h7fb7e90ff7839cc4;
    assign coff[4793] = 64'h544f63d29fb063d9;
    assign coff[4794] = 64'hf7839cc4804816f1;
    assign coff[4795] = 64'h9fb063d9abb09c2e;
    assign coff[4796] = 64'h604f9c27abb09c2e;
    assign coff[4797] = 64'h087c633c804816f1;
    assign coff[4798] = 64'habb09c2e9fb063d9;
    assign coff[4799] = 64'h804816f1f7839cc4;
    assign coff[4800] = 64'h618782fdad1a30d9;
    assign coff[4801] = 64'h0a589c94806b37cf;
    assign coff[4802] = 64'had1a30d99e787d03;
    assign coff[4803] = 64'h806b37cff5a7636c;
    assign coff[4804] = 64'h7f94c831f5a7636c;
    assign coff[4805] = 64'h52e5cf279e787d03;
    assign coff[4806] = 64'hf5a7636c806b37cf;
    assign coff[4807] = 64'h9e787d03ad1a30d9;
    assign coff[4808] = 64'h79d43532d8bc4207;
    assign coff[4809] = 64'h3a61bcfd8e16f3a9;
    assign coff[4810] = 64'hd8bc4207862bcace;
    assign coff[4811] = 64'h8e16f3a9c59e4303;
    assign coff[4812] = 64'h71e90c57c59e4303;
    assign coff[4813] = 64'h2743bdf9862bcace;
    assign coff[4814] = 64'hc59e43038e16f3a9;
    assign coff[4815] = 64'h862bcaced8bc4207;
    assign coff[4816] = 64'h6fd3f001c1b8e1bf;
    assign coff[4817] = 64'h2309859384e38118;
    assign coff[4818] = 64'hc1b8e1bf902c0fff;
    assign coff[4819] = 64'h84e38118dcf67a6d;
    assign coff[4820] = 64'h7b1c7ee8dcf67a6d;
    assign coff[4821] = 64'h3e471e41902c0fff;
    assign coff[4822] = 64'hdcf67a6d84e38118;
    assign coff[4823] = 64'h902c0fffc1b8e1bf;
    assign coff[4824] = 64'h7f25eec7f141eab5;
    assign coff[4825] = 64'h4f7b992d9bab0ac3;
    assign coff[4826] = 64'hf141eab580da1139;
    assign coff[4827] = 64'h9bab0ac3b08466d3;
    assign coff[4828] = 64'h6454f53db08466d3;
    assign coff[4829] = 64'h0ebe154b80da1139;
    assign coff[4830] = 64'hb08466d39bab0ac3;
    assign coff[4831] = 64'h80da1139f141eab5;
    assign coff[4832] = 64'h692f6328b70f9fac;
    assign coff[4833] = 64'h16cd2c9f820c1912;
    assign coff[4834] = 64'hb70f9fac96d09cd8;
    assign coff[4835] = 64'h820c1912e932d361;
    assign coff[4836] = 64'h7df3e6eee932d361;
    assign coff[4837] = 64'h48f0605496d09cd8;
    assign coff[4838] = 64'he932d361820c1912;
    assign coff[4839] = 64'h96d09cd8b70f9fac;
    assign coff[4840] = 64'h7d174564e4dda385;
    assign coff[4841] = 64'h45440d90945c4f09;
    assign coff[4842] = 64'he4dda38582e8ba9c;
    assign coff[4843] = 64'h945c4f09babbf270;
    assign coff[4844] = 64'h6ba3b0f7babbf270;
    assign coff[4845] = 64'h1b225c7b82e8ba9c;
    assign coff[4846] = 64'hbabbf270945c4f09;
    assign coff[4847] = 64'h82e8ba9ce4dda385;
    assign coff[4848] = 64'h7564c8f8ccfbae4d;
    assign coff[4849] = 64'h2eef7ce588ea6e83;
    assign coff[4850] = 64'hccfbae4d8a9b3708;
    assign coff[4851] = 64'h88ea6e83d110831b;
    assign coff[4852] = 64'h7715917dd110831b;
    assign coff[4853] = 64'h330451b38a9b3708;
    assign coff[4854] = 64'hd110831b88ea6e83;
    assign coff[4855] = 64'h8a9b3708ccfbae4d;
    assign coff[4856] = 64'h7ffb1ee9fdca8a99;
    assign coff[4857] = 64'h58ef2f6ba3f122b2;
    assign coff[4858] = 64'hfdca8a998004e117;
    assign coff[4859] = 64'ha3f122b2a710d095;
    assign coff[4860] = 64'h5c0edd4ea710d095;
    assign coff[4861] = 64'h023575678004e117;
    assign coff[4862] = 64'ha710d095a3f122b2;
    assign coff[4863] = 64'h8004e117fdca8a99;
    assign coff[4864] = 64'h5c43304da7471a07;
    assign coff[4865] = 64'h0280d81380064460;
    assign coff[4866] = 64'ha7471a07a3bccfb3;
    assign coff[4867] = 64'h80064460fd7f27ed;
    assign coff[4868] = 64'h7ff9bba0fd7f27ed;
    assign coff[4869] = 64'h58b8e5f9a3bccfb3;
    assign coff[4870] = 64'hfd7f27ed80064460;
    assign coff[4871] = 64'ha3bccfb3a7471a07;
    assign coff[4872] = 64'h77312287d156b0b7;
    assign coff[4873] = 64'h33496f628ab9588e;
    assign coff[4874] = 64'hd156b0b788cedd79;
    assign coff[4875] = 64'h8ab9588eccb6909e;
    assign coff[4876] = 64'h7546a772ccb6909e;
    assign coff[4877] = 64'h2ea94f4988cedd79;
    assign coff[4878] = 64'hccb6909e8ab9588e;
    assign coff[4879] = 64'h88cedd79d156b0b7;
    assign coff[4880] = 64'h6bcc6b53bafb6615;
    assign coff[4881] = 64'h1b6c070582f8cc0d;
    assign coff[4882] = 64'hbafb6615943394ad;
    assign coff[4883] = 64'h82f8cc0de493f8fb;
    assign coff[4884] = 64'h7d0733f3e493f8fb;
    assign coff[4885] = 64'h450499eb943394ad;
    assign coff[4886] = 64'he493f8fb82f8cc0d;
    assign coff[4887] = 64'h943394adbafb6615;
    assign coff[4888] = 64'h7e013f74e97d088c;
    assign coff[4889] = 64'h492e493396fba605;
    assign coff[4890] = 64'he97d088c81fec08c;
    assign coff[4891] = 64'h96fba605b6d1b6cd;
    assign coff[4892] = 64'h690459fbb6d1b6cd;
    assign coff[4893] = 64'h1682f77481fec08c;
    assign coff[4894] = 64'hb6d1b6cd96fba605;
    assign coff[4895] = 64'h81fec08ce97d088c;
    assign coff[4896] = 64'h6483b58cb0bf8e4a;
    assign coff[4897] = 64'h0f08f83680e2d666;
    assign coff[4898] = 64'hb0bf8e4a9b7c4a74;
    assign coff[4899] = 64'h80e2d666f0f707ca;
    assign coff[4900] = 64'h7f1d299af0f707ca;
    assign coff[4901] = 64'h4f4071b69b7c4a74;
    assign coff[4902] = 64'hf0f707ca80e2d666;
    assign coff[4903] = 64'h9b7c4a74b0bf8e4a;
    assign coff[4904] = 64'h7b310d07dd3f053c;
    assign coff[4905] = 64'h3e88f2ae9050d2a9;
    assign coff[4906] = 64'hdd3f053c84cef2f9;
    assign coff[4907] = 64'h9050d2a9c1770d52;
    assign coff[4908] = 64'h6faf2d57c1770d52;
    assign coff[4909] = 64'h22c0fac484cef2f9;
    assign coff[4910] = 64'hc1770d529050d2a9;
    assign coff[4911] = 64'h84cef2f9dd3f053c;
    assign coff[4912] = 64'h720b5c57c5e16667;
    assign coff[4913] = 64'h278b7a84864300e7;
    assign coff[4914] = 64'hc5e166678df4a3a9;
    assign coff[4915] = 64'h864300e7d874857c;
    assign coff[4916] = 64'h79bcff19d874857c;
    assign coff[4917] = 64'h3a1e99998df4a3a9;
    assign coff[4918] = 64'hd874857c864300e7;
    assign coff[4919] = 64'h8df4a3a9c5e16667;
    assign coff[4920] = 64'h7f9aca37f5f28bfd;
    assign coff[4921] = 64'h531f33d59ea96299;
    assign coff[4922] = 64'hf5f28bfd806535c9;
    assign coff[4923] = 64'h9ea96299ace0cc2b;
    assign coff[4924] = 64'h61569d67ace0cc2b;
    assign coff[4925] = 64'h0a0d7403806535c9;
    assign coff[4926] = 64'hace0cc2b9ea96299;
    assign coff[4927] = 64'h806535c9f5f28bfd;
    assign coff[4928] = 64'h60813519abe96625;
    assign coff[4929] = 64'h08c79d3a804d2cbd;
    assign coff[4930] = 64'habe966259f7ecae7;
    assign coff[4931] = 64'h804d2cbdf73862c6;
    assign coff[4932] = 64'h7fb2d343f73862c6;
    assign coff[4933] = 64'h541699db9f7ecae7;
    assign coff[4934] = 64'hf73862c6804d2cbd;
    assign coff[4935] = 64'h9f7ecae7abe96625;
    assign coff[4936] = 64'h79568250d73e499a;
    assign coff[4937] = 64'h38fac30e8d61bd89;
    assign coff[4938] = 64'hd73e499a86a97db0;
    assign coff[4939] = 64'h8d61bd89c7053cf2;
    assign coff[4940] = 64'h729e4277c7053cf2;
    assign coff[4941] = 64'h28c1b66686a97db0;
    assign coff[4942] = 64'hc7053cf28d61bd89;
    assign coff[4943] = 64'h86a97db0d73e499a;
    assign coff[4944] = 64'h6f0e22a3c05ac603;
    assign coff[4945] = 64'h2186172b8477cebd;
    assign coff[4946] = 64'hc05ac60390f1dd5d;
    assign coff[4947] = 64'h8477cebdde79e8d5;
    assign coff[4948] = 64'h7b883143de79e8d5;
    assign coff[4949] = 64'h3fa539fd90f1dd5d;
    assign coff[4950] = 64'hde79e8d58477cebd;
    assign coff[4951] = 64'h90f1dd5dc05ac603;
    assign coff[4952] = 64'h7ef52b00efb2c365;
    assign coff[4953] = 64'h4e3edf4d9ab3479d;
    assign coff[4954] = 64'hefb2c365810ad500;
    assign coff[4955] = 64'h9ab3479db1c120b3;
    assign coff[4956] = 64'h654cb863b1c120b3;
    assign coff[4957] = 64'h104d3c9b810ad500;
    assign coff[4958] = 64'hb1c120b39ab3479d;
    assign coff[4959] = 64'h810ad500efb2c365;
    assign coff[4960] = 64'h68483891b5c696da;
    assign coff[4961] = 64'h15410d7081c6e50d;
    assign coff[4962] = 64'hb5c696da97b7c76f;
    assign coff[4963] = 64'h81c6e50deabef290;
    assign coff[4964] = 64'h7e391af3eabef290;
    assign coff[4965] = 64'h4a39692697b7c76f;
    assign coff[4966] = 64'heabef29081c6e50d;
    assign coff[4967] = 64'h97b7c76fb5c696da;
    assign coff[4968] = 64'h7cbf9e03e3552fdf;
    assign coff[4969] = 64'h43f0912b9384c8b8;
    assign coff[4970] = 64'he3552fdf834061fd;
    assign coff[4971] = 64'h9384c8b8bc0f6ed5;
    assign coff[4972] = 64'h6c7b3748bc0f6ed5;
    assign coff[4973] = 64'h1caad021834061fd;
    assign coff[4974] = 64'hbc0f6ed59384c8b8;
    assign coff[4975] = 64'h834061fde3552fdf;
    assign coff[4976] = 64'h74c2407dcb8bded1;
    assign coff[4977] = 64'h2d787a7288594757;
    assign coff[4978] = 64'hcb8bded18b3dbf83;
    assign coff[4979] = 64'h88594757d287858e;
    assign coff[4980] = 64'h77a6b8a9d287858e;
    assign coff[4981] = 64'h3474212f8b3dbf83;
    assign coff[4982] = 64'hd287858e88594757;
    assign coff[4983] = 64'h8b3dbf83cb8bded1;
    assign coff[4984] = 64'h7ff1b6f6fc3887b3;
    assign coff[4985] = 64'h57cc44eca2db858e;
    assign coff[4986] = 64'hfc3887b3800e490a;
    assign coff[4987] = 64'ha2db858ea833bb14;
    assign coff[4988] = 64'h5d247a72a833bb14;
    assign coff[4989] = 64'h03c7784d800e490a;
    assign coff[4990] = 64'ha833bb14a2db858e;
    assign coff[4991] = 64'h800e490afc3887b3;
    assign coff[4992] = 64'h5e697a39a9919616;
    assign coff[4993] = 64'h05a4aa09801fdc86;
    assign coff[4994] = 64'ha9919616a19685c7;
    assign coff[4995] = 64'h801fdc86fa5b55f7;
    assign coff[4996] = 64'h7fe0237afa5b55f7;
    assign coff[4997] = 64'h566e69eaa19685c7;
    assign coff[4998] = 64'hfa5b55f7801fdc86;
    assign coff[4999] = 64'ha19685c7a9919616;
    assign coff[5000] = 64'h784d18f4d4471e29;
    assign coff[5001] = 64'h362646098c0499c4;
    assign coff[5002] = 64'hd4471e2987b2e70c;
    assign coff[5003] = 64'h8c0499c4c9d9b9f7;
    assign coff[5004] = 64'h73fb663cc9d9b9f7;
    assign coff[5005] = 64'h2bb8e1d787b2e70c;
    assign coff[5006] = 64'hc9d9b9f78c0499c4;
    assign coff[5007] = 64'h87b2e70cd4471e29;
    assign coff[5008] = 64'h6d75b786bda5f862;
    assign coff[5009] = 64'h1e7b68c283aeb797;
    assign coff[5010] = 64'hbda5f862928a487a;
    assign coff[5011] = 64'h83aeb797e184973e;
    assign coff[5012] = 64'h7c514869e184973e;
    assign coff[5013] = 64'h425a079e928a487a;
    assign coff[5014] = 64'he184973e83aeb797;
    assign coff[5015] = 64'h928a487abda5f862;
    assign coff[5016] = 64'h7e84f67eec9666cd;
    assign coff[5017] = 64'h4bbc6b2598cf820b;
    assign coff[5018] = 64'hec9666cd817b0982;
    assign coff[5019] = 64'h98cf820bb44394db;
    assign coff[5020] = 64'h67307df5b44394db;
    assign coff[5021] = 64'h13699933817b0982;
    assign coff[5022] = 64'hb44394db98cf820b;
    assign coff[5023] = 64'h817b0982ec9666cd;
    assign coff[5024] = 64'h666ddcd3b33d2771;
    assign coff[5025] = 64'h12266913814b18c3;
    assign coff[5026] = 64'hb33d27719992232d;
    assign coff[5027] = 64'h814b18c3edd996ed;
    assign coff[5028] = 64'h7eb4e73dedd996ed;
    assign coff[5029] = 64'h4cc2d88f9992232d;
    assign coff[5030] = 64'hedd996ed814b18c3;
    assign coff[5031] = 64'h9992232db33d2771;
    assign coff[5032] = 64'h7c01e534e047a875;
    assign coff[5033] = 64'h4141c9fb91e25032;
    assign coff[5034] = 64'he047a87583fe1acc;
    assign coff[5035] = 64'h91e25032bebe3605;
    assign coff[5036] = 64'h6e1dafcebebe3605;
    assign coff[5037] = 64'h1fb8578b83fe1acc;
    assign coff[5038] = 64'hbebe360591e25032;
    assign coff[5039] = 64'h83fe1acce047a875;
    assign coff[5040] = 64'h736fb4ecc8b25f06;
    assign coff[5041] = 64'h2a8541c38744d51b;
    assign coff[5042] = 64'hc8b25f068c904b14;
    assign coff[5043] = 64'h8744d51bd57abe3d;
    assign coff[5044] = 64'h78bb2ae5d57abe3d;
    assign coff[5045] = 64'h374da0fa8c904b14;
    assign coff[5046] = 64'hd57abe3d8744d51b;
    assign coff[5047] = 64'h8c904b14c8b25f06;
    assign coff[5048] = 64'h7fd01b63f915014c;
    assign coff[5049] = 64'h557c53b6a0bb1ba2;
    assign coff[5050] = 64'hf915014c802fe49d;
    assign coff[5051] = 64'ha0bb1ba2aa83ac4a;
    assign coff[5052] = 64'h5f44e45eaa83ac4a;
    assign coff[5053] = 64'h06eafeb4802fe49d;
    assign coff[5054] = 64'haa83ac4aa0bb1ba2;
    assign coff[5055] = 64'h802fe49df915014c;
    assign coff[5056] = 64'h628a0e50ae4e2db6;
    assign coff[5057] = 64'h0be935d2808e2e0a;
    assign coff[5058] = 64'hae4e2db69d75f1b0;
    assign coff[5059] = 64'h808e2e0af416ca2e;
    assign coff[5060] = 64'h7f71d1f6f416ca2e;
    assign coff[5061] = 64'h51b1d24a9d75f1b0;
    assign coff[5062] = 64'hf416ca2e808e2e0a;
    assign coff[5063] = 64'h9d75f1b0ae4e2db6;
    assign coff[5064] = 64'h7a4d35b0da3bbdf9;
    assign coff[5065] = 64'h3bc676b98ed08e05;
    assign coff[5066] = 64'hda3bbdf985b2ca50;
    assign coff[5067] = 64'h8ed08e05c4398947;
    assign coff[5068] = 64'h712f71fbc4398947;
    assign coff[5069] = 64'h25c4420785b2ca50;
    assign coff[5070] = 64'hc43989478ed08e05;
    assign coff[5071] = 64'h85b2ca50da3bbdf9;
    assign coff[5072] = 64'h70956db1c3196422;
    assign coff[5073] = 64'h248b9a2f8553f27e;
    assign coff[5074] = 64'hc31964228f6a924f;
    assign coff[5075] = 64'h8553f27edb7465d1;
    assign coff[5076] = 64'h7aac0d82db7465d1;
    assign coff[5077] = 64'h3ce69bde8f6a924f;
    assign coff[5078] = 64'hdb7465d18553f27e;
    assign coff[5079] = 64'h8f6a924fc3196422;
    assign coff[5080] = 64'h7f51cbabf2d1a385;
    assign coff[5081] = 64'h50b5429a9ca6ac23;
    assign coff[5082] = 64'hf2d1a38580ae3455;
    assign coff[5083] = 64'h9ca6ac23af4abd66;
    assign coff[5084] = 64'h635953ddaf4abd66;
    assign coff[5085] = 64'h0d2e5c7b80ae3455;
    assign coff[5086] = 64'haf4abd669ca6ac23;
    assign coff[5087] = 64'h80ae3455f2d1a385;
    assign coff[5088] = 64'h6a127f9fb85b785e;
    assign coff[5089] = 64'h18586ac38256282e;
    assign coff[5090] = 64'hb85b785e95ed8061;
    assign coff[5091] = 64'h8256282ee7a7953d;
    assign coff[5092] = 64'h7da9d7d2e7a7953d;
    assign coff[5093] = 64'h47a487a295ed8061;
    assign coff[5094] = 64'he7a7953d8256282e;
    assign coff[5095] = 64'h95ed8061b85b785e;
    assign coff[5096] = 64'h7d6a1a31e66722f7;
    assign coff[5097] = 64'h4694de569537fbb2;
    assign coff[5098] = 64'he66722f78295e5cf;
    assign coff[5099] = 64'h9537fbb2b96b21aa;
    assign coff[5100] = 64'h6ac8044eb96b21aa;
    assign coff[5101] = 64'h1998dd098295e5cf;
    assign coff[5102] = 64'hb96b21aa9537fbb2;
    assign coff[5103] = 64'h8295e5cfe66722f7;
    assign coff[5104] = 64'h7602cad5ce6d754c;
    assign coff[5105] = 64'h3064b01d89802cfc;
    assign coff[5106] = 64'hce6d754c89fd352b;
    assign coff[5107] = 64'h89802cfccf9b4fe3;
    assign coff[5108] = 64'h767fd304cf9b4fe3;
    assign coff[5109] = 64'h31928ab489fd352b;
    assign coff[5110] = 64'hcf9b4fe389802cfc;
    assign coff[5111] = 64'h89fd352bce6d754c;
    assign coff[5112] = 64'h7fff97c1ff5ca34b;
    assign coff[5113] = 64'h5a0eac2ea50a4c68;
    assign coff[5114] = 64'hff5ca34b8000683f;
    assign coff[5115] = 64'ha50a4c68a5f153d2;
    assign coff[5116] = 64'h5af5b398a5f153d2;
    assign coff[5117] = 64'h00a35cb58000683f;
    assign coff[5118] = 64'ha5f153d2a50a4c68;
    assign coff[5119] = 64'h8000683fff5ca34b;
    assign coff[5120] = 64'h5ae40311a5df796b;
    assign coff[5121] = 64'h008a3acb80004aa4;
    assign coff[5122] = 64'ha5df796ba51bfcef;
    assign coff[5123] = 64'h80004aa4ff75c535;
    assign coff[5124] = 64'h7fffb55cff75c535;
    assign coff[5125] = 64'h5a208695a51bfcef;
    assign coff[5126] = 64'hff75c53580004aa4;
    assign coff[5127] = 64'ha51bfcefa5df796b;
    assign coff[5128] = 64'h76765038cf840c65;
    assign coff[5129] = 64'h317b5de089f37ba9;
    assign coff[5130] = 64'hcf840c658989afc8;
    assign coff[5131] = 64'h89f37ba9ce84a220;
    assign coff[5132] = 64'h760c8457ce84a220;
    assign coff[5133] = 64'h307bf39b8989afc8;
    assign coff[5134] = 64'hce84a22089f37ba9;
    assign coff[5135] = 64'h8989afc8cf840c65;
    assign coff[5136] = 64'h6aba266eb9562b9c;
    assign coff[5137] = 64'h19803c868290e194;
    assign coff[5138] = 64'hb9562b9c9545d992;
    assign coff[5139] = 64'h8290e194e67fc37a;
    assign coff[5140] = 64'h7d6f1e6ce67fc37a;
    assign coff[5141] = 64'h46a9d4649545d992;
    assign coff[5142] = 64'he67fc37a8290e194;
    assign coff[5143] = 64'h9545d992b9562b9c;
    assign coff[5144] = 64'h7da50dabe78ee92c;
    assign coff[5145] = 64'h478fb27b95df7145;
    assign coff[5146] = 64'he78ee92c825af255;
    assign coff[5147] = 64'h95df7145b8704d85;
    assign coff[5148] = 64'h6a208ebbb8704d85;
    assign coff[5149] = 64'h187116d4825af255;
    assign coff[5150] = 64'hb8704d8595df7145;
    assign coff[5151] = 64'h825af255e78ee92c;
    assign coff[5152] = 64'h6349791faf373d22;
    assign coff[5153] = 64'h0d155c7380aba03b;
    assign coff[5154] = 64'haf373d229cb686e1;
    assign coff[5155] = 64'h80aba03bf2eaa38d;
    assign coff[5156] = 64'h7f545fc5f2eaa38d;
    assign coff[5157] = 64'h50c8c2de9cb686e1;
    assign coff[5158] = 64'hf2eaa38d80aba03b;
    assign coff[5159] = 64'h9cb686e1af373d22;
    assign coff[5160] = 64'h7aa4de2ddb5c505a;
    assign coff[5161] = 64'h3cd07f9f8f5e9f46;
    assign coff[5162] = 64'hdb5c505a855b21d3;
    assign coff[5163] = 64'h8f5e9f46c32f8061;
    assign coff[5164] = 64'h70a160bac32f8061;
    assign coff[5165] = 64'h24a3afa6855b21d3;
    assign coff[5166] = 64'hc32f80618f5e9f46;
    assign coff[5167] = 64'h855b21d3db5c505a;
    assign coff[5168] = 64'h7123b32bc423511d;
    assign coff[5169] = 64'h25ac3dc085ab6250;
    assign coff[5170] = 64'hc423511d8edc4cd5;
    assign coff[5171] = 64'h85ab6250da53c240;
    assign coff[5172] = 64'h7a549db0da53c240;
    assign coff[5173] = 64'h3bdcaee38edc4cd5;
    assign coff[5174] = 64'hda53c24085ab6250;
    assign coff[5175] = 64'h8edc4cd5c423511d;
    assign coff[5176] = 64'h7f6f78cbf3fdc459;
    assign coff[5177] = 64'h519e77979d65e92b;
    assign coff[5178] = 64'hf3fdc45980908735;
    assign coff[5179] = 64'h9d65e92bae618869;
    assign coff[5180] = 64'h629a16d5ae618869;
    assign coff[5181] = 64'h0c023ba780908735;
    assign coff[5182] = 64'hae6188699d65e92b;
    assign coff[5183] = 64'h80908735f3fdc459;
    assign coff[5184] = 64'h5f34198eaa70f930;
    assign coff[5185] = 64'h06d1e5fe802e8b58;
    assign coff[5186] = 64'haa70f930a0cbe672;
    assign coff[5187] = 64'h802e8b58f92e1a02;
    assign coff[5188] = 64'h7fd174a8f92e1a02;
    assign coff[5189] = 64'h558f06d0a0cbe672;
    assign coff[5190] = 64'hf92e1a02802e8b58;
    assign coff[5191] = 64'ha0cbe672aa70f930;
    assign coff[5192] = 64'h78b2cf41d5630a74;
    assign coff[5193] = 64'h3736f5738c857176;
    assign coff[5194] = 64'hd5630a74874d30bf;
    assign coff[5195] = 64'h8c857176c8c90a8d;
    assign coff[5196] = 64'h737a8e8ac8c90a8d;
    assign coff[5197] = 64'h2a9cf58c874d30bf;
    assign coff[5198] = 64'hc8c90a8d8c857176;
    assign coff[5199] = 64'h874d30bfd5630a74;
    assign coff[5200] = 64'h6e10dd82bea8983f;
    assign coff[5201] = 64'h1f9ffda483f7e2c3;
    assign coff[5202] = 64'hbea8983f91ef227e;
    assign coff[5203] = 64'h83f7e2c3e060025c;
    assign coff[5204] = 64'h7c081d3de060025c;
    assign coff[5205] = 64'h415767c191ef227e;
    assign coff[5206] = 64'he060025c83f7e2c3;
    assign coff[5207] = 64'h91ef227ebea8983f;
    assign coff[5208] = 64'h7eb1547aedc0b64e;
    assign coff[5209] = 64'h4caeba6e998312b7;
    assign coff[5210] = 64'hedc0b64e814eab86;
    assign coff[5211] = 64'h998312b7b3514592;
    assign coff[5212] = 64'h667ced49b3514592;
    assign coff[5213] = 64'h123f49b2814eab86;
    assign coff[5214] = 64'hb3514592998312b7;
    assign coff[5215] = 64'h814eab86edc0b64e;
    assign coff[5216] = 64'h67219d10b42f5373;
    assign coff[5217] = 64'h1350c14481773c2b;
    assign coff[5218] = 64'hb42f537398de62f0;
    assign coff[5219] = 64'h81773c2becaf3ebc;
    assign coff[5220] = 64'h7e88c3d5ecaf3ebc;
    assign coff[5221] = 64'h4bd0ac8d98de62f0;
    assign coff[5222] = 64'hecaf3ebc81773c2b;
    assign coff[5223] = 64'h98de62f0b42f5373;
    assign coff[5224] = 64'h7c4b49d2e16c2ef4;
    assign coff[5225] = 64'h42448849927d4363;
    assign coff[5226] = 64'he16c2ef483b4b62e;
    assign coff[5227] = 64'h927d4363bdbb77b7;
    assign coff[5228] = 64'h6d82bc9dbdbb77b7;
    assign coff[5229] = 64'h1e93d10c83b4b62e;
    assign coff[5230] = 64'hbdbb77b7927d4363;
    assign coff[5231] = 64'h83b4b62ee16c2ef4;
    assign coff[5232] = 64'h73f0c226c9c2f51e;
    assign coff[5233] = 64'h2ba1420087aa53a6;
    assign coff[5234] = 64'hc9c2f51e8c0f3dda;
    assign coff[5235] = 64'h87aa53a6d45ebe00;
    assign coff[5236] = 64'h7855ac5ad45ebe00;
    assign coff[5237] = 64'h363d0ae28c0f3dda;
    assign coff[5238] = 64'hd45ebe0087aa53a6;
    assign coff[5239] = 64'h8c0f3ddac9c2f51e;
    assign coff[5240] = 64'h7fdf055afa423a59;
    assign coff[5241] = 64'h565bde95a1858f16;
    assign coff[5242] = 64'hfa423a598020faa6;
    assign coff[5243] = 64'ha1858f16a9a4216b;
    assign coff[5244] = 64'h5e7a70eaa9a4216b;
    assign coff[5245] = 64'h05bdc5a78020faa6;
    assign coff[5246] = 64'ha9a4216ba1858f16;
    assign coff[5247] = 64'h8020faa6fa423a59;
    assign coff[5248] = 64'h5d133b72a82172eb;
    assign coff[5249] = 64'h03ae590d800d8d8b;
    assign coff[5250] = 64'ha82172eba2ecc48e;
    assign coff[5251] = 64'h800d8d8bfc51a6f3;
    assign coff[5252] = 64'h7ff27275fc51a6f3;
    assign coff[5253] = 64'h57de8d15a2ecc48e;
    assign coff[5254] = 64'hfc51a6f3800d8d8b;
    assign coff[5255] = 64'ha2ecc48ea82172eb;
    assign coff[5256] = 64'h779dc8c0d270081b;
    assign coff[5257] = 64'h345d333c8b337528;
    assign coff[5258] = 64'hd270081b88623740;
    assign coff[5259] = 64'h8b337528cba2ccc4;
    assign coff[5260] = 64'h74cc8ad8cba2ccc4;
    assign coff[5261] = 64'h2d8ff7e588623740;
    assign coff[5262] = 64'hcba2ccc48b337528;
    assign coff[5263] = 64'h88623740d270081b;
    assign coff[5264] = 64'h6c6dde2bbbfa2347;
    assign coff[5265] = 64'h1c925109833ac36c;
    assign coff[5266] = 64'hbbfa2347939221d5;
    assign coff[5267] = 64'h833ac36ce36daef7;
    assign coff[5268] = 64'h7cc53c94e36daef7;
    assign coff[5269] = 64'h4405dcb9939221d5;
    assign coff[5270] = 64'he36daef7833ac36c;
    assign coff[5271] = 64'h939221d5bbfa2347;
    assign coff[5272] = 64'h7e34ec2beaa62a4f;
    assign coff[5273] = 64'h4a24edee97a93687;
    assign coff[5274] = 64'heaa62a4f81cb13d5;
    assign coff[5275] = 64'h97a93687b5db1212;
    assign coff[5276] = 64'h6856c979b5db1212;
    assign coff[5277] = 64'h1559d5b181cb13d5;
    assign coff[5278] = 64'hb5db121297a93687;
    assign coff[5279] = 64'h81cb13d5eaa62a4f;
    assign coff[5280] = 64'h653d5962b1ad3e55;
    assign coff[5281] = 64'h10344eb48107a409;
    assign coff[5282] = 64'hb1ad3e559ac2a69e;
    assign coff[5283] = 64'h8107a409efcbb14c;
    assign coff[5284] = 64'h7ef85bf7efcbb14c;
    assign coff[5285] = 64'h4e52c1ab9ac2a69e;
    assign coff[5286] = 64'hefcbb14c8107a409;
    assign coff[5287] = 64'h9ac2a69eb1ad3e55;
    assign coff[5288] = 64'h7b8199cade61a815;
    assign coff[5289] = 64'h3f8f6a8590e56056;
    assign coff[5290] = 64'hde61a815847e6636;
    assign coff[5291] = 64'h90e56056c070957b;
    assign coff[5292] = 64'h6f1a9faac070957b;
    assign coff[5293] = 64'h219e57eb847e6636;
    assign coff[5294] = 64'hc070957b90e56056;
    assign coff[5295] = 64'h847e6636de61a815;
    assign coff[5296] = 64'h72931027c6eebcb5;
    assign coff[5297] = 64'h28a9e28186a17f5f;
    assign coff[5298] = 64'hc6eebcb58d6cefd9;
    assign coff[5299] = 64'h86a17f5fd7561d7f;
    assign coff[5300] = 64'h795e80a1d7561d7f;
    assign coff[5301] = 64'h3911434b8d6cefd9;
    assign coff[5302] = 64'hd7561d7f86a17f5f;
    assign coff[5303] = 64'h8d6cefd9c6eebcb5;
    assign coff[5304] = 64'h7fb1177bf71f501e;
    assign coff[5305] = 64'h5403a5619f6e4a06;
    assign coff[5306] = 64'hf71f501e804ee885;
    assign coff[5307] = 64'h9f6e4a06abfc5a9f;
    assign coff[5308] = 64'h6091b5faabfc5a9f;
    assign coff[5309] = 64'h08e0afe2804ee885;
    assign coff[5310] = 64'habfc5a9f9f6e4a06;
    assign coff[5311] = 64'h804ee885f71f501e;
    assign coff[5312] = 64'h6146495daccdb103;
    assign coff[5313] = 64'h09f465b580633ef3;
    assign coff[5314] = 64'haccdb1039eb9b6a3;
    assign coff[5315] = 64'h80633ef3f60b9a4b;
    assign coff[5316] = 64'h7f9cc10df60b9a4b;
    assign coff[5317] = 64'h53324efd9eb9b6a3;
    assign coff[5318] = 64'hf60b9a4b80633ef3;
    assign coff[5319] = 64'h9eb9b6a3accdb103;
    assign coff[5320] = 64'h79b53903d85c9f04;
    assign coff[5321] = 64'h3a0833fc8de93c74;
    assign coff[5322] = 64'hd85c9f04864ac6fd;
    assign coff[5323] = 64'h8de93c74c5f7cc04;
    assign coff[5324] = 64'h7216c38cc5f7cc04;
    assign coff[5325] = 64'h27a360fc864ac6fd;
    assign coff[5326] = 64'hc5f7cc048de93c74;
    assign coff[5327] = 64'h864ac6fdd85c9f04;
    assign coff[5328] = 64'h6fa2e3d7c16120a9;
    assign coff[5329] = 64'h22a8c9cf84c8226e;
    assign coff[5330] = 64'hc16120a9905d1c29;
    assign coff[5331] = 64'h84c8226edd573631;
    assign coff[5332] = 64'h7b37dd92dd573631;
    assign coff[5333] = 64'h3e9edf57905d1c29;
    assign coff[5334] = 64'hdd57363184c8226e;
    assign coff[5335] = 64'h905d1c29c16120a9;
    assign coff[5336] = 64'h7f1a3368f0de12a3;
    assign coff[5337] = 64'h4f2cb3c79b6cbcc4;
    assign coff[5338] = 64'hf0de12a380e5cc98;
    assign coff[5339] = 64'h9b6cbcc4b0d34c39;
    assign coff[5340] = 64'h6493433cb0d34c39;
    assign coff[5341] = 64'h0f21ed5d80e5cc98;
    assign coff[5342] = 64'hb0d34c399b6cbcc4;
    assign coff[5343] = 64'h80e5cc98f0de12a3;
    assign coff[5344] = 64'h68f5f97db6bd197c;
    assign coff[5345] = 64'h166a395381fa576c;
    assign coff[5346] = 64'hb6bd197c970a0683;
    assign coff[5347] = 64'h81fa576ce995c6ad;
    assign coff[5348] = 64'h7e05a894e995c6ad;
    assign coff[5349] = 64'h4942e684970a0683;
    assign coff[5350] = 64'he995c6ad81fa576c;
    assign coff[5351] = 64'h970a0683b6bd197c;
    assign coff[5352] = 64'h7d01cf29e47b6ce9;
    assign coff[5353] = 64'h44ef6e0b94260989;
    assign coff[5354] = 64'he47b6ce982fe30d7;
    assign coff[5355] = 64'h94260989bb1091f5;
    assign coff[5356] = 64'h6bd9f677bb1091f5;
    assign coff[5357] = 64'h1b84931782fe30d7;
    assign coff[5358] = 64'hbb1091f594260989;
    assign coff[5359] = 64'h82fe30d7e47b6ce9;
    assign coff[5360] = 64'h753c933acc9f8aac;
    assign coff[5361] = 64'h2e91e72588c5b650;
    assign coff[5362] = 64'hcc9f8aac8ac36cc6;
    assign coff[5363] = 64'h88c5b650d16e18db;
    assign coff[5364] = 64'h773a49b0d16e18db;
    assign coff[5365] = 64'h336075548ac36cc6;
    assign coff[5366] = 64'hd16e18db88c5b650;
    assign coff[5367] = 64'h8ac36cc6cc9f8aac;
    assign coff[5368] = 64'h7ff93b54fd660739;
    assign coff[5369] = 64'h58a6c6a5a3ab65d0;
    assign coff[5370] = 64'hfd6607398006c4ac;
    assign coff[5371] = 64'ha3ab65d0a759395b;
    assign coff[5372] = 64'h5c549a30a759395b;
    assign coff[5373] = 64'h0299f8c78006c4ac;
    assign coff[5374] = 64'ha759395ba3ab65d0;
    assign coff[5375] = 64'h8006c4acfd660739;
    assign coff[5376] = 64'h5bfd6534a6febef4;
    assign coff[5377] = 64'h021c545780047488;
    assign coff[5378] = 64'ha6febef4a4029acc;
    assign coff[5379] = 64'h80047488fde3aba9;
    assign coff[5380] = 64'h7ffb8b78fde3aba9;
    assign coff[5381] = 64'h5901410ca4029acc;
    assign coff[5382] = 64'hfde3aba980047488;
    assign coff[5383] = 64'ha4029acca6febef4;
    assign coff[5384] = 64'h770c57f5d0f9222f;
    assign coff[5385] = 64'h32ed43de8a9134e8;
    assign coff[5386] = 64'hd0f9222f88f3a80b;
    assign coff[5387] = 64'h8a9134e8cd12bc22;
    assign coff[5388] = 64'h756ecb18cd12bc22;
    assign coff[5389] = 64'h2f06ddd188f3a80b;
    assign coff[5390] = 64'hcd12bc228a9134e8;
    assign coff[5391] = 64'h88f3a80bd0f9222f;
    assign coff[5392] = 64'h6b961536baa6d13a;
    assign coff[5393] = 64'h1b09cc3482e3691b;
    assign coff[5394] = 64'hbaa6d13a9469eaca;
    assign coff[5395] = 64'h82e3691be4f633cc;
    assign coff[5396] = 64'h7d1c96e5e4f633cc;
    assign coff[5397] = 64'h45592ec69469eaca;
    assign coff[5398] = 64'he4f633cc82e3691b;
    assign coff[5399] = 64'h9469eacabaa6d13a;
    assign coff[5400] = 64'h7def6a60e91a18bf;
    assign coff[5401] = 64'h48dbb7be96c24c8f;
    assign coff[5402] = 64'he91a18bf821095a0;
    assign coff[5403] = 64'h96c24c8fb7244842;
    assign coff[5404] = 64'h693db371b7244842;
    assign coff[5405] = 64'h16e5e741821095a0;
    assign coff[5406] = 64'hb724484296c24c8f;
    assign coff[5407] = 64'h821095a0e91a18bf;
    assign coff[5408] = 64'h64455810b070b520;
    assign coff[5409] = 64'h0ea51dd880d72ea3;
    assign coff[5410] = 64'hb070b5209bbaa7f0;
    assign coff[5411] = 64'h80d72ea3f15ae228;
    assign coff[5412] = 64'h7f28d15df15ae228;
    assign coff[5413] = 64'h4f8f4ae09bbaa7f0;
    assign coff[5414] = 64'hf15ae22880d72ea3;
    assign coff[5415] = 64'h9bbaa7f0b070b520;
    assign coff[5416] = 64'h7b159b5fdcde4eda;
    assign coff[5417] = 64'h3e3127f9901fd7ba;
    assign coff[5418] = 64'hdcde4eda84ea64a1;
    assign coff[5419] = 64'h901fd7bac1ced807;
    assign coff[5420] = 64'h6fe02846c1ced807;
    assign coff[5421] = 64'h2321b12684ea64a1;
    assign coff[5422] = 64'hc1ced807901fd7ba;
    assign coff[5423] = 64'h84ea64a1dcde4eda;
    assign coff[5424] = 64'h71dd938fc587e661;
    assign coff[5425] = 64'h272bd16d86241780;
    assign coff[5426] = 64'hc587e6618e226c71;
    assign coff[5427] = 64'h86241780d8d42e93;
    assign coff[5428] = 64'h79dbe880d8d42e93;
    assign coff[5429] = 64'h3a78199f8e226c71;
    assign coff[5430] = 64'hd8d42e9386241780;
    assign coff[5431] = 64'h8e226c71c587e661;
    assign coff[5432] = 64'h7f92bdadf58e56b1;
    assign coff[5433] = 64'h52d2a7329e683800;
    assign coff[5434] = 64'hf58e56b1806d4253;
    assign coff[5435] = 64'h9e683800ad2d58ce;
    assign coff[5436] = 64'h6197c800ad2d58ce;
    assign coff[5437] = 64'h0a71a94f806d4253;
    assign coff[5438] = 64'had2d58ce9e683800;
    assign coff[5439] = 64'h806d4253f58e56b1;
    assign coff[5440] = 64'h603f0c69ab9db4b0;
    assign coff[5441] = 64'h08634f3e80466edb;
    assign coff[5442] = 64'hab9db4b09fc0f397;
    assign coff[5443] = 64'h80466edbf79cb0c2;
    assign coff[5444] = 64'h7fb99125f79cb0c2;
    assign coff[5445] = 64'h54624b509fc0f397;
    assign coff[5446] = 64'hf79cb0c280466edb;
    assign coff[5447] = 64'h9fc0f397ab9db4b0;
    assign coff[5448] = 64'h79365a49d6df09c6;
    assign coff[5449] = 64'h38a0ac298d35207d;
    assign coff[5450] = 64'hd6df09c686c9a5b7;
    assign coff[5451] = 64'h8d35207dc75f53d7;
    assign coff[5452] = 64'h72cadf83c75f53d7;
    assign coff[5453] = 64'h2920f63a86c9a5b7;
    assign coff[5454] = 64'hc75f53d78d35207d;
    assign coff[5455] = 64'h86c9a5b7d6df09c6;
    assign coff[5456] = 64'h6edc03bcc003a0b3;
    assign coff[5457] = 64'h21250749845da07e;
    assign coff[5458] = 64'hc003a0b39123fc44;
    assign coff[5459] = 64'h845da07ededaf8b7;
    assign coff[5460] = 64'h7ba25f82dedaf8b7;
    assign coff[5461] = 64'h3ffc5f4d9123fc44;
    assign coff[5462] = 64'hdedaf8b7845da07e;
    assign coff[5463] = 64'h9123fc44c003a0b3;
    assign coff[5464] = 64'h7ee83632ef4f121b;
    assign coff[5465] = 64'h4def37b09a75f2ac;
    assign coff[5466] = 64'hef4f121b8117c9ce;
    assign coff[5467] = 64'h9a75f2acb210c850;
    assign coff[5468] = 64'h658a0d54b210c850;
    assign coff[5469] = 64'h10b0ede58117c9ce;
    assign coff[5470] = 64'hb210c8509a75f2ac;
    assign coff[5471] = 64'h8117c9ceef4f121b;
    assign coff[5472] = 64'h680dccc1b574c69d;
    assign coff[5473] = 64'h14dde44581b65a99;
    assign coff[5474] = 64'hb574c69d97f2333f;
    assign coff[5475] = 64'h81b65a99eb221bbb;
    assign coff[5476] = 64'h7e49a567eb221bbb;
    assign coff[5477] = 64'h4a8b396397f2333f;
    assign coff[5478] = 64'heb221bbb81b65a99;
    assign coff[5479] = 64'h97f2333fb574c69d;
    assign coff[5480] = 64'h7ca8f3a7e2f33e94;
    assign coff[5481] = 64'h439b48c9934f8e1c;
    assign coff[5482] = 64'he2f33e9483570c59;
    assign coff[5483] = 64'h934f8e1cbc64b737;
    assign coff[5484] = 64'h6cb071e4bc64b737;
    assign coff[5485] = 64'h1d0cc16c83570c59;
    assign coff[5486] = 64'hbc64b737934f8e1c;
    assign coff[5487] = 64'h83570c59e2f33e94;
    assign coff[5488] = 64'h7498ea11cb303b49;
    assign coff[5489] = 64'h2d1a73258835b5d9;
    assign coff[5490] = 64'hcb303b498b6715ef;
    assign coff[5491] = 64'h8835b5d9d2e58cdb;
    assign coff[5492] = 64'h77ca4a27d2e58cdb;
    assign coff[5493] = 64'h34cfc4b78b6715ef;
    assign coff[5494] = 64'hd2e58cdb8835b5d9;
    assign coff[5495] = 64'h8b6715efcb303b49;
    assign coff[5496] = 64'h7fee97a7fbd40c33;
    assign coff[5497] = 64'h57830276a296ad7d;
    assign coff[5498] = 64'hfbd40c3380116859;
    assign coff[5499] = 64'ha296ad7da87cfd8a;
    assign coff[5500] = 64'h5d695283a87cfd8a;
    assign coff[5501] = 64'h042bf3cd80116859;
    assign coff[5502] = 64'ha87cfd8aa296ad7d;
    assign coff[5503] = 64'h80116859fbd40c33;
    assign coff[5504] = 64'h5e257b17a9478a1c;
    assign coff[5505] = 64'h0540396f801b9554;
    assign coff[5506] = 64'ha9478a1ca1da84e9;
    assign coff[5507] = 64'h801b9554fabfc691;
    assign coff[5508] = 64'h7fe46aacfabfc691;
    assign coff[5509] = 64'h56b875e4a1da84e9;
    assign coff[5510] = 64'hfabfc691801b9554;
    assign coff[5511] = 64'ha1da84e9a9478a1c;
    assign coff[5512] = 64'h782a9cfed3e8afb3;
    assign coff[5513] = 64'h35cb1dcc8bda3626;
    assign coff[5514] = 64'hd3e8afb387d56302;
    assign coff[5515] = 64'h8bda3626ca34e234;
    assign coff[5516] = 64'h7425c9daca34e234;
    assign coff[5517] = 64'h2c17504d87d56302;
    assign coff[5518] = 64'hca34e2348bda3626;
    assign coff[5519] = 64'h87d56302d3e8afb3;
    assign coff[5520] = 64'h6d4178fdbd5014ad;
    assign coff[5521] = 64'h1e19bbe08396ed29;
    assign coff[5522] = 64'hbd5014ad92be8703;
    assign coff[5523] = 64'h8396ed29e1e64420;
    assign coff[5524] = 64'h7c6912d7e1e64420;
    assign coff[5525] = 64'h42afeb5392be8703;
    assign coff[5526] = 64'he1e644208396ed29;
    assign coff[5527] = 64'h92be8703bd5014ad;
    assign coff[5528] = 64'h7e75905dec330e99;
    assign coff[5529] = 64'h4b6b485a98942643;
    assign coff[5530] = 64'hec330e99818a6fa3;
    assign coff[5531] = 64'h98942643b494b7a6;
    assign coff[5532] = 64'h676bd9bdb494b7a6;
    assign coff[5533] = 64'h13ccf167818a6fa3;
    assign coff[5534] = 64'hb494b7a698942643;
    assign coff[5535] = 64'h818a6fa3ec330e99;
    assign coff[5536] = 64'h66317385b2eccc8c;
    assign coff[5537] = 64'h11c2dfa2813cfe91;
    assign coff[5538] = 64'hb2eccc8c99ce8c7b;
    assign coff[5539] = 64'h813cfe91ee3d205e;
    assign coff[5540] = 64'h7ec3016fee3d205e;
    assign coff[5541] = 64'h4d13337499ce8c7b;
    assign coff[5542] = 64'hee3d205e813cfe91;
    assign coff[5543] = 64'h99ce8c7bb2eccc8c;
    assign coff[5544] = 64'h7be8d544dfe64d1c;
    assign coff[5545] = 64'h40eb39c391af317c;
    assign coff[5546] = 64'hdfe64d1c84172abc;
    assign coff[5547] = 64'h91af317cbf14c63d;
    assign coff[5548] = 64'h6e50ce84bf14c63d;
    assign coff[5549] = 64'h2019b2e484172abc;
    assign coff[5550] = 64'hbf14c63d91af317c;
    assign coff[5551] = 64'h84172abcdfe64d1c;
    assign coff[5552] = 64'h734421f6c857c642;
    assign coff[5553] = 64'h2a26624087239518;
    assign coff[5554] = 64'hc857c6428cbbde0a;
    assign coff[5555] = 64'h87239518d5d99dc0;
    assign coff[5556] = 64'h78dc6ae8d5d99dc0;
    assign coff[5557] = 64'h37a839be8cbbde0a;
    assign coff[5558] = 64'hd5d99dc087239518;
    assign coff[5559] = 64'h8cbbde0ac857c642;
    assign coff[5560] = 64'h7fca8508f8b0a129;
    assign coff[5561] = 64'h55316663a0781522;
    assign coff[5562] = 64'hf8b0a12980357af8;
    assign coff[5563] = 64'ha0781522aace999d;
    assign coff[5564] = 64'h5f87eadeaace999d;
    assign coff[5565] = 64'h074f5ed780357af8;
    assign coff[5566] = 64'haace999da0781522;
    assign coff[5567] = 64'h80357af8f8b0a129;
    assign coff[5568] = 64'h6249c645ae00e271;
    assign coff[5569] = 64'h0b8519ed8084fa82;
    assign coff[5570] = 64'hae00e2719db639bb;
    assign coff[5571] = 64'h8084fa82f47ae613;
    assign coff[5572] = 64'h7f7b057ef47ae613;
    assign coff[5573] = 64'h51ff1d8f9db639bb;
    assign coff[5574] = 64'hf47ae6138084fa82;
    assign coff[5575] = 64'h9db639bbae00e271;
    assign coff[5576] = 64'h7a2f668cd9dbbb77;
    assign coff[5577] = 64'h3b6d7f108ea1be6c;
    assign coff[5578] = 64'hd9dbbb7785d09974;
    assign coff[5579] = 64'h8ea1be6cc49280f0;
    assign coff[5580] = 64'h715e4194c49280f0;
    assign coff[5581] = 64'h2624448985d09974;
    assign coff[5582] = 64'hc49280f08ea1be6c;
    assign coff[5583] = 64'h85d09974d9dbbb77;
    assign coff[5584] = 64'h70657626c2c10aa7;
    assign coff[5585] = 64'h242b364485376477;
    assign coff[5586] = 64'hc2c10aa78f9a89da;
    assign coff[5587] = 64'h85376477dbd4c9bc;
    assign coff[5588] = 64'h7ac89b89dbd4c9bc;
    assign coff[5589] = 64'h3d3ef5598f9a89da;
    assign coff[5590] = 64'hdbd4c9bc85376477;
    assign coff[5591] = 64'h8f9a89dac2c10aa7;
    assign coff[5592] = 64'h7f474a30f26da885;
    assign coff[5593] = 64'h506722739c67677c;
    assign coff[5594] = 64'hf26da88580b8b5d0;
    assign coff[5595] = 64'h9c67677caf98dd8d;
    assign coff[5596] = 64'h63989884af98dd8d;
    assign coff[5597] = 64'h0d92577b80b8b5d0;
    assign coff[5598] = 64'haf98dd8d9c67677c;
    assign coff[5599] = 64'h80b8b5d0f26da885;
    assign coff[5600] = 64'h69da1a50b8083f67;
    assign coff[5601] = 64'h17f5b12982433004;
    assign coff[5602] = 64'hb8083f679625e5b0;
    assign coff[5603] = 64'h82433004e80a4ed7;
    assign coff[5604] = 64'h7dbccffce80a4ed7;
    assign coff[5605] = 64'h47f7c0999625e5b0;
    assign coff[5606] = 64'he80a4ed782433004;
    assign coff[5607] = 64'h9625e5b0b8083f67;
    assign coff[5608] = 64'h7d55d8e9e604aad4;
    assign coff[5609] = 64'h4640eaf29500ad66;
    assign coff[5610] = 64'he604aad482aa2717;
    assign coff[5611] = 64'h9500ad66b9bf150e;
    assign coff[5612] = 64'h6aff529ab9bf150e;
    assign coff[5613] = 64'h19fb552c82aa2717;
    assign coff[5614] = 64'hb9bf150e9500ad66;
    assign coff[5615] = 64'h82aa2717e604aad4;
    assign coff[5616] = 64'h75dbb753ce10d51f;
    assign coff[5617] = 64'h30078f86895a4f7e;
    assign coff[5618] = 64'hce10d51f8a2448ad;
    assign coff[5619] = 64'h895a4f7ecff8707a;
    assign coff[5620] = 64'h76a5b082cff8707a;
    assign coff[5621] = 64'h31ef2ae18a2448ad;
    assign coff[5622] = 64'hcff8707a895a4f7e;
    assign coff[5623] = 64'h8a2448adce10d51f;
    assign coff[5624] = 64'h7ffeeff8fef81bec;
    assign coff[5625] = 64'h59c71fe3a4c3ad64;
    assign coff[5626] = 64'hfef81bec80011008;
    assign coff[5627] = 64'ha4c3ad64a638e01d;
    assign coff[5628] = 64'h5b3c529ca638e01d;
    assign coff[5629] = 64'h0107e41480011008;
    assign coff[5630] = 64'ha638e01da4c3ad64;
    assign coff[5631] = 64'h80011008fef81bec;
    assign coff[5632] = 64'h5b7124f2a66eadb0;
    assign coff[5633] = 64'h015349348001c1ae;
    assign coff[5634] = 64'ha66eadb0a48edb0e;
    assign coff[5635] = 64'h8001c1aefeacb6cc;
    assign coff[5636] = 64'h7ffe3e52feacb6cc;
    assign coff[5637] = 64'h59915250a48edb0e;
    assign coff[5638] = 64'hfeacb6cc8001c1ae;
    assign coff[5639] = 64'ha48edb0ea66eadb0;
    assign coff[5640] = 64'h76c1e699d03e5c60;
    assign coff[5641] = 64'h32348ecf8a41c706;
    assign coff[5642] = 64'hd03e5c60893e1967;
    assign coff[5643] = 64'h8a41c706cdcb7131;
    assign coff[5644] = 64'h75be38facdcb7131;
    assign coff[5645] = 64'h2fc1a3a0893e1967;
    assign coff[5646] = 64'hcdcb71318a41c706;
    assign coff[5647] = 64'h893e1967d03e5c60;
    assign coff[5648] = 64'h6b28a206b9fe280d;
    assign coff[5649] = 64'h1a4524c682b98aca;
    assign coff[5650] = 64'hb9fe280d94d75dfa;
    assign coff[5651] = 64'h82b98acae5badb3a;
    assign coff[5652] = 64'h7d467536e5badb3a;
    assign coff[5653] = 64'h4601d7f394d75dfa;
    assign coff[5654] = 64'he5badb3a82b98aca;
    assign coff[5655] = 64'h94d75dfab9fe280d;
    assign coff[5656] = 64'h7dcad736e85463c2;
    assign coff[5657] = 64'h48360e3296505c88;
    assign coff[5658] = 64'he85463c2823528ca;
    assign coff[5659] = 64'h96505c88b7c9f1ce;
    assign coff[5660] = 64'h69afa378b7c9f1ce;
    assign coff[5661] = 64'h17ab9c3e823528ca;
    assign coff[5662] = 64'hb7c9f1ce96505c88;
    assign coff[5663] = 64'h823528cae85463c2;
    assign coff[5664] = 64'h63c7e3b1afd39638;
    assign coff[5665] = 64'h0ddd4e4080c0ca73;
    assign coff[5666] = 64'hafd396389c381c4f;
    assign coff[5667] = 64'h80c0ca73f222b1c0;
    assign coff[5668] = 64'h7f3f358df222b1c0;
    assign coff[5669] = 64'h502c69c89c381c4f;
    assign coff[5670] = 64'hf222b1c080c0ca73;
    assign coff[5671] = 64'h9c381c4fafd39638;
    assign coff[5672] = 64'h7addd45bdc1d2354;
    assign coff[5673] = 64'h3d811fac8fbeb103;
    assign coff[5674] = 64'hdc1d235485222ba5;
    assign coff[5675] = 64'h8fbeb103c27ee054;
    assign coff[5676] = 64'h70414efdc27ee054;
    assign coff[5677] = 64'h23e2dcac85222ba5;
    assign coff[5678] = 64'hc27ee0548fbeb103;
    assign coff[5679] = 64'h85222ba5dc1d2354;
    assign coff[5680] = 64'h71812f65c4d552c1;
    assign coff[5681] = 64'h266c36fe85e72647;
    assign coff[5682] = 64'hc4d552c18e7ed09b;
    assign coff[5683] = 64'h85e72647d993c902;
    assign coff[5684] = 64'h7a18d9b9d993c902;
    assign coff[5685] = 64'h3b2aad3f8e7ed09b;
    assign coff[5686] = 64'hd993c90285e72647;
    assign coff[5687] = 64'h8e7ed09bc4d552c1;
    assign coff[5688] = 64'h7f81b88af4c5ffab;
    assign coff[5689] = 64'h5238f4d49de6978f;
    assign coff[5690] = 64'hf4c5ffab807e4776;
    assign coff[5691] = 64'h9de6978fadc70b2c;
    assign coff[5692] = 64'h62196871adc70b2c;
    assign coff[5693] = 64'h0b3a0055807e4776;
    assign coff[5694] = 64'hadc70b2c9de6978f;
    assign coff[5695] = 64'h807e4776f4c5ffab;
    assign coff[5696] = 64'h5fba0914ab06ee1b;
    assign coff[5697] = 64'h079aa4008039df77;
    assign coff[5698] = 64'hab06ee1ba045f6ec;
    assign coff[5699] = 64'h8039df77f8655c00;
    assign coff[5700] = 64'h7fc62089f8655c00;
    assign coff[5701] = 64'h54f911e5a045f6ec;
    assign coff[5702] = 64'hf8655c008039df77;
    assign coff[5703] = 64'ha045f6ecab06ee1b;
    assign coff[5704] = 64'h78f529fed620d675;
    assign coff[5705] = 64'h37ec15cb8cdcbaee;
    assign coff[5706] = 64'hd620d675870ad602;
    assign coff[5707] = 64'h8cdcbaeec813ea35;
    assign coff[5708] = 64'h73234512c813ea35;
    assign coff[5709] = 64'h29df298b870ad602;
    assign coff[5710] = 64'hc813ea358cdcbaee;
    assign coff[5711] = 64'h870ad602d620d675;
    assign coff[5712] = 64'h6e76f8e7bf55ccb2;
    assign coff[5713] = 64'h2062aa6b842a28da;
    assign coff[5714] = 64'hbf55ccb291890719;
    assign coff[5715] = 64'h842a28dadf9d5595;
    assign coff[5716] = 64'h7bd5d726df9d5595;
    assign coff[5717] = 64'h40aa334e91890719;
    assign coff[5718] = 64'hdf9d5595842a28da;
    assign coff[5719] = 64'h91890719bf55ccb2;
    assign coff[5720] = 64'h7ecd61c5ee87cea7;
    assign coff[5721] = 64'h4d4f587099fc04d6;
    assign coff[5722] = 64'hee87cea781329e3b;
    assign coff[5723] = 64'h99fc04d6b2b0a790;
    assign coff[5724] = 64'h6603fb2ab2b0a790;
    assign coff[5725] = 64'h1178315981329e3b;
    assign coff[5726] = 64'hb2b0a79099fc04d6;
    assign coff[5727] = 64'h81329e3bee87cea7;
    assign coff[5728] = 64'h679834b6b4d1b048;
    assign coff[5729] = 64'h14176b8e81962f6d;
    assign coff[5730] = 64'hb4d1b0489867cb4a;
    assign coff[5731] = 64'h81962f6debe89472;
    assign coff[5732] = 64'h7e69d093ebe89472;
    assign coff[5733] = 64'h4b2e4fb89867cb4a;
    assign coff[5734] = 64'hebe8947281962f6d;
    assign coff[5735] = 64'h9867cb4ab4d1b048;
    assign coff[5736] = 64'h7c7ab84ee22f91fc;
    assign coff[5737] = 64'h42f03b1e92e5e226;
    assign coff[5738] = 64'he22f91fc838547b2;
    assign coff[5739] = 64'h92e5e226bd0fc4e2;
    assign coff[5740] = 64'h6d1a1ddabd0fc4e2;
    assign coff[5741] = 64'h1dd06e04838547b2;
    assign coff[5742] = 64'hbd0fc4e292e5e226;
    assign coff[5743] = 64'h838547b2e22f91fc;
    assign coff[5744] = 64'h7445658dca79562b;
    assign coff[5745] = 64'h2c5e114f87ef70a0;
    assign coff[5746] = 64'hca79562b8bba9a73;
    assign coff[5747] = 64'h87ef70a0d3a1eeb1;
    assign coff[5748] = 64'h78108f60d3a1eeb1;
    assign coff[5749] = 64'h3586a9d58bba9a73;
    assign coff[5750] = 64'hd3a1eeb187ef70a0;
    assign coff[5751] = 64'h8bba9a73ca79562b;
    assign coff[5752] = 64'h7fe76c4cfb0b1d28;
    assign coff[5753] = 64'h56efdbc7a20daa62;
    assign coff[5754] = 64'hfb0b1d28801893b4;
    assign coff[5755] = 64'ha20daa62a9102439;
    assign coff[5756] = 64'h5df2559ea9102439;
    assign coff[5757] = 64'h04f4e2d8801893b4;
    assign coff[5758] = 64'ha9102439a20daa62;
    assign coff[5759] = 64'h801893b4fb0b1d28;
    assign coff[5760] = 64'h5d9ccec2a8b412d1;
    assign coff[5761] = 64'h04774ec18013f39e;
    assign coff[5762] = 64'ha8b412d1a263313e;
    assign coff[5763] = 64'h8013f39efb88b13f;
    assign coff[5764] = 64'h7fec0c62fb88b13f;
    assign coff[5765] = 64'h574bed2fa263313e;
    assign coff[5766] = 64'hfb88b13f8013f39e;
    assign coff[5767] = 64'ha263313ea8b412d1;
    assign coff[5768] = 64'h77e4c6c9d32c2499;
    assign coff[5769] = 64'h35146a008b8645f5;
    assign coff[5770] = 64'hd32c2499881b3937;
    assign coff[5771] = 64'h8b8645f5caeb9600;
    assign coff[5772] = 64'h7479ba0bcaeb9600;
    assign coff[5773] = 64'h2cd3db67881b3937;
    assign coff[5774] = 64'hcaeb96008b8645f5;
    assign coff[5775] = 64'h881b3937d32c2499;
    assign coff[5776] = 64'h6cd831dcbca4c8e1;
    assign coff[5777] = 64'h1d562aa683683e95;
    assign coff[5778] = 64'hbca4c8e19327ce24;
    assign coff[5779] = 64'h83683e95e2a9d55a;
    assign coff[5780] = 64'h7c97c16be2a9d55a;
    assign coff[5781] = 64'h435b371f9327ce24;
    assign coff[5782] = 64'he2a9d55a83683e95;
    assign coff[5783] = 64'h9327ce24bca4c8e1;
    assign coff[5784] = 64'h7e55da20eb6c8312;
    assign coff[5785] = 64'h4ac87767981e2e3c;
    assign coff[5786] = 64'heb6c831281aa25e0;
    assign coff[5787] = 64'h981e2e3cb5378899;
    assign coff[5788] = 64'h67e1d1c4b5378899;
    assign coff[5789] = 64'h14937cee81aa25e0;
    assign coff[5790] = 64'hb5378899981e2e3c;
    assign coff[5791] = 64'h81aa25e0eb6c8312;
    assign coff[5792] = 64'h65b7e3f1b24ca594;
    assign coff[5793] = 64'h10fbac1e8121b4c8;
    assign coff[5794] = 64'hb24ca5949a481c0f;
    assign coff[5795] = 64'h8121b4c8ef0453e2;
    assign coff[5796] = 64'h7ede4b38ef0453e2;
    assign coff[5797] = 64'h4db35a6c9a481c0f;
    assign coff[5798] = 64'hef0453e28121b4c8;
    assign coff[5799] = 64'h9a481c0fb24ca594;
    assign coff[5800] = 64'h7bb5d026df23d20e;
    assign coff[5801] = 64'h403da1659149c053;
    assign coff[5802] = 64'hdf23d20e844a2fda;
    assign coff[5803] = 64'h9149c053bfc25e9b;
    assign coff[5804] = 64'h6eb63fadbfc25e9b;
    assign coff[5805] = 64'h20dc2df2844a2fda;
    assign coff[5806] = 64'hbfc25e9b9149c053;
    assign coff[5807] = 64'h844a2fdadf23d20e;
    assign coff[5808] = 64'h72ec26d6c7a2fbf3;
    assign coff[5809] = 64'h2968557686e1f4cf;
    assign coff[5810] = 64'hc7a2fbf38d13d92a;
    assign coff[5811] = 64'h86e1f4cfd697aa8a;
    assign coff[5812] = 64'h791e0b31d697aa8a;
    assign coff[5813] = 64'h385d040d8d13d92a;
    assign coff[5814] = 64'hd697aa8a86e1f4cf;
    assign coff[5815] = 64'h8d13d92ac7a2fbf3;
    assign coff[5816] = 64'h7fbe6bdbf7e7eea7;
    assign coff[5817] = 64'h549aee429ff2b914;
    assign coff[5818] = 64'hf7e7eea780419425;
    assign coff[5819] = 64'h9ff2b914ab6511be;
    assign coff[5820] = 64'h600d46ecab6511be;
    assign coff[5821] = 64'h0818115980419425;
    assign coff[5822] = 64'hab6511be9ff2b914;
    assign coff[5823] = 64'h80419425f7e7eea7;
    assign coff[5824] = 64'h61c88074ad66e3d3;
    assign coff[5825] = 64'h0abccd1180737f5f;
    assign coff[5826] = 64'had66e3d39e377f8c;
    assign coff[5827] = 64'h80737f5ff54332ef;
    assign coff[5828] = 64'h7f8c80a1f54332ef;
    assign coff[5829] = 64'h52991c2d9e377f8c;
    assign coff[5830] = 64'hf54332ef80737f5f;
    assign coff[5831] = 64'h9e377f8cad66e3d3;
    assign coff[5832] = 64'h79f2e63ad91bfd43;
    assign coff[5833] = 64'h3abb21fb8e44f121;
    assign coff[5834] = 64'hd91bfd43860d19c6;
    assign coff[5835] = 64'h8e44f121c544de05;
    assign coff[5836] = 64'h71bb0edfc544de05;
    assign coff[5837] = 64'h26e402bd860d19c6;
    assign coff[5838] = 64'hc544de058e44f121;
    assign coff[5839] = 64'h860d19c6d91bfd43;
    assign coff[5840] = 64'h7004b731c210c940;
    assign coff[5841] = 64'h236a2bba84ff2bb3;
    assign coff[5842] = 64'hc210c9408ffb48cf;
    assign coff[5843] = 64'h84ff2bb3dc95d446;
    assign coff[5844] = 64'h7b00d44ddc95d446;
    assign coff[5845] = 64'h3def36c08ffb48cf;
    assign coff[5846] = 64'hdc95d44684ff2bb3;
    assign coff[5847] = 64'h8ffb48cfc210c940;
    assign coff[5848] = 64'h7f315bb7f1a5cbdf;
    assign coff[5849] = 64'h4fca4d8d9be996a6;
    assign coff[5850] = 64'hf1a5cbdf80cea449;
    assign coff[5851] = 64'h9be996a6b035b273;
    assign coff[5852] = 64'h6416695ab035b273;
    assign coff[5853] = 64'h0e5a342180cea449;
    assign coff[5854] = 64'hb035b2739be996a6;
    assign coff[5855] = 64'h80cea449f1a5cbdf;
    assign coff[5856] = 64'h69688bf1b76252db;
    assign coff[5857] = 64'h173011d9821e286b;
    assign coff[5858] = 64'hb76252db9697740f;
    assign coff[5859] = 64'h821e286be8cfee27;
    assign coff[5860] = 64'h7de1d795e8cfee27;
    assign coff[5861] = 64'h489dad259697740f;
    assign coff[5862] = 64'he8cfee27821e286b;
    assign coff[5863] = 64'h9697740fb76252db;
    assign coff[5864] = 64'h7d2c6e76e53feade;
    assign coff[5865] = 64'h4598825a9492d6ef;
    assign coff[5866] = 64'he53feade82d3918a;
    assign coff[5867] = 64'h9492d6efba677da6;
    assign coff[5868] = 64'h6b6d2911ba677da6;
    assign coff[5869] = 64'h1ac0152282d3918a;
    assign coff[5870] = 64'hba677da69492d6ef;
    assign coff[5871] = 64'h82d3918ae53feade;
    assign coff[5872] = 64'h758cb64ccd57f167;
    assign coff[5873] = 64'h2f4cf5b0890f702b;
    assign coff[5874] = 64'hcd57f1678a7349b4;
    assign coff[5875] = 64'h890f702bd0b30a50;
    assign coff[5876] = 64'h76f08fd5d0b30a50;
    assign coff[5877] = 64'h32a80e998a7349b4;
    assign coff[5878] = 64'hd0b30a50890f702b;
    assign coff[5879] = 64'h8a7349b4cd57f167;
    assign coff[5880] = 64'h7ffcb38cfe2f0f55;
    assign coff[5881] = 64'h59376155a437185e;
    assign coff[5882] = 64'hfe2f0f5580034c74;
    assign coff[5883] = 64'ha437185ea6c89eab;
    assign coff[5884] = 64'h5bc8e7a2a6c89eab;
    assign coff[5885] = 64'h01d0f0ab80034c74;
    assign coff[5886] = 64'ha6c89eaba437185e;
    assign coff[5887] = 64'h80034c74fe2f0f55;
    assign coff[5888] = 64'h5c88c27ca78fabd4;
    assign coff[5889] = 64'h02e55a448008632a;
    assign coff[5890] = 64'ha78fabd4a3773d84;
    assign coff[5891] = 64'h8008632afd1aa5bc;
    assign coff[5892] = 64'h7ff79cd6fd1aa5bc;
    assign coff[5893] = 64'h5870542ca3773d84;
    assign coff[5894] = 64'hfd1aa5bc8008632a;
    assign coff[5895] = 64'ha3773d84a78fabd4;
    assign coff[5896] = 64'h7755a394d1b45c08;
    assign coff[5897] = 64'h33a57b448ae1c48b;
    assign coff[5898] = 64'hd1b45c0888aa5c6c;
    assign coff[5899] = 64'h8ae1c48bcc5a84bc;
    assign coff[5900] = 64'h751e3b75cc5a84bc;
    assign coff[5901] = 64'h2e4ba3f888aa5c6c;
    assign coff[5902] = 64'hcc5a84bc8ae1c48b;
    assign coff[5903] = 64'h88aa5c6cd1b45c08;
    assign coff[5904] = 64'h6c027ef1bb502583;
    assign coff[5905] = 64'h1bce30ec830e7c1f;
    assign coff[5906] = 64'hbb50258393fd810f;
    assign coff[5907] = 64'h830e7c1fe431cf14;
    assign coff[5908] = 64'h7cf183e1e431cf14;
    assign coff[5909] = 64'h44afda7d93fd810f;
    assign coff[5910] = 64'he431cf14830e7c1f;
    assign coff[5911] = 64'h93fd810fbb502583;
    assign coff[5912] = 64'h7e12c6cee9e0063c;
    assign coff[5913] = 64'h4980ad8497354043;
    assign coff[5914] = 64'he9e0063c81ed3932;
    assign coff[5915] = 64'h97354043b67f527c;
    assign coff[5916] = 64'h68cabfbdb67f527c;
    assign coff[5917] = 64'h161ff9c481ed3932;
    assign coff[5918] = 64'hb67f527c97354043;
    assign coff[5919] = 64'h81ed3932e9e0063c;
    assign coff[5920] = 64'h64c1d507b10e9856;
    assign coff[5921] = 64'h0f6cc94e80eecc93;
    assign coff[5922] = 64'hb10e98569b3e2af9;
    assign coff[5923] = 64'h80eecc93f09336b2;
    assign coff[5924] = 64'h7f11336df09336b2;
    assign coff[5925] = 64'h4ef167aa9b3e2af9;
    assign coff[5926] = 64'hf09336b280eecc93;
    assign coff[5927] = 64'h9b3e2af9b10e9856;
    assign coff[5928] = 64'h7b4c32b1dd9fd10f;
    assign coff[5929] = 64'h3ee096d19082127c;
    assign coff[5930] = 64'hdd9fd10f84b3cd4f;
    assign coff[5931] = 64'h9082127cc11f692f;
    assign coff[5932] = 64'h6f7ded84c11f692f;
    assign coff[5933] = 64'h22602ef184b3cd4f;
    assign coff[5934] = 64'hc11f692f9082127c;
    assign coff[5935] = 64'h84b3cd4fdd9fd10f;
    assign coff[5936] = 64'h7238dec5c63b0a46;
    assign coff[5937] = 64'h27eb0b3686623566;
    assign coff[5938] = 64'hc63b0a468dc7213b;
    assign coff[5939] = 64'h86623566d814f4ca;
    assign coff[5940] = 64'h799dca9ad814f4ca;
    assign coff[5941] = 64'h39c4f5ba8dc7213b;
    assign coff[5942] = 64'hd814f4ca86623566;
    assign coff[5943] = 64'h8dc7213bc63b0a46;
    assign coff[5944] = 64'h7fa2880bf656c77c;
    assign coff[5945] = 64'h536b8d339eeac93e;
    assign coff[5946] = 64'hf656c77c805d77f5;
    assign coff[5947] = 64'h9eeac93eac9472cd;
    assign coff[5948] = 64'h611536c2ac9472cd;
    assign coff[5949] = 64'h09a93884805d77f5;
    assign coff[5950] = 64'hac9472cd9eeac93e;
    assign coff[5951] = 64'h805d77f5f656c77c;
    assign coff[5952] = 64'h60c32243ac354b7a;
    assign coff[5953] = 64'h092be5ca80543965;
    assign coff[5954] = 64'hac354b7a9f3cddbd;
    assign coff[5955] = 64'h80543965f6d41a36;
    assign coff[5956] = 64'h7fabc69bf6d41a36;
    assign coff[5957] = 64'h53cab4869f3cddbd;
    assign coff[5958] = 64'hf6d41a3680543965;
    assign coff[5959] = 64'h9f3cddbdac354b7a;
    assign coff[5960] = 64'h79765f7fd79da293;
    assign coff[5961] = 64'h3954b6cd8d8ea148;
    assign coff[5962] = 64'hd79da2938689a081;
    assign coff[5963] = 64'h8d8ea148c6ab4933;
    assign coff[5964] = 64'h72715eb8c6ab4933;
    assign coff[5965] = 64'h28625d6d8689a081;
    assign coff[5966] = 64'hc6ab49338d8ea148;
    assign coff[5967] = 64'h8689a081d79da293;
    assign coff[5968] = 64'h6f3ffd09c0b21295;
    assign coff[5969] = 64'h21e7126084924930;
    assign coff[5970] = 64'hc0b2129590c002f7;
    assign coff[5971] = 64'h84924930de18eda0;
    assign coff[5972] = 64'h7b6db6d0de18eda0;
    assign coff[5973] = 64'h3f4ded6b90c002f7;
    assign coff[5974] = 64'hde18eda084924930;
    assign coff[5975] = 64'h90c002f7c0b21295;
    assign coff[5976] = 64'h7f01d17df0167ebd;
    assign coff[5977] = 64'h4e8e56a59af0db0b;
    assign coff[5978] = 64'hf0167ebd80fe2e83;
    assign coff[5979] = 64'h9af0db0bb171a95b;
    assign coff[5980] = 64'h650f24f5b171a95b;
    assign coff[5981] = 64'h0fe9814380fe2e83;
    assign coff[5982] = 64'hb171a95b9af0db0b;
    assign coff[5983] = 64'h80fe2e83f0167ebd;
    assign coff[5984] = 64'h6882640eb61894df;
    assign coff[5985] = 64'h15a4297f81d7bd5e;
    assign coff[5986] = 64'hb61894df977d9bf2;
    assign coff[5987] = 64'h81d7bd5eea5bd681;
    assign coff[5988] = 64'h7e2842a2ea5bd681;
    assign coff[5989] = 64'h49e76b21977d9bf2;
    assign coff[5990] = 64'hea5bd68181d7bd5e;
    assign coff[5991] = 64'h977d9bf2b61894df;
    assign coff[5992] = 64'h7cd5fb6ae3b732d9;
    assign coff[5993] = 64'h4445afa493ba463f;
    assign coff[5994] = 64'he3b732d9832a0496;
    assign coff[5995] = 64'h93ba463fbbba505c;
    assign coff[5996] = 64'h6c45b9c1bbba505c;
    assign coff[5997] = 64'h1c48cd27832a0496;
    assign coff[5998] = 64'hbbba505c93ba463f;
    assign coff[5999] = 64'h832a0496e3b732d9;
    assign coff[6000] = 64'h74eb4ee3cbe7a2b5;
    assign coff[6001] = 64'h2dd665b2887d22a4;
    assign coff[6002] = 64'hcbe7a2b58b14b11d;
    assign coff[6003] = 64'h887d22a4d2299a4e;
    assign coff[6004] = 64'h7782dd5cd2299a4e;
    assign coff[6005] = 64'h34185d4b8b14b11d;
    assign coff[6006] = 64'hd2299a4e887d22a4;
    assign coff[6007] = 64'h8b14b11dcbe7a2b5;
    assign coff[6008] = 64'h7ff48759fc9d0588;
    assign coff[6009] = 64'h58155139a3209713;
    assign coff[6010] = 64'hfc9d0588800b78a7;
    assign coff[6011] = 64'ha3209713a7eaaec7;
    assign coff[6012] = 64'h5cdf68eda7eaaec7;
    assign coff[6013] = 64'h0362fa78800b78a7;
    assign coff[6014] = 64'ha7eaaec7a3209713;
    assign coff[6015] = 64'h800b78a7fc9d0588;
    assign coff[6016] = 64'h5ead3f1fa9dbd761;
    assign coff[6017] = 64'h0609172980247299;
    assign coff[6018] = 64'ha9dbd761a152c0e1;
    assign coff[6019] = 64'h80247299f9f6e8d7;
    assign coff[6020] = 64'h7fdb8d67f9f6e8d7;
    assign coff[6021] = 64'h5624289fa152c0e1;
    assign coff[6022] = 64'hf9f6e8d780247299;
    assign coff[6023] = 64'ha152c0e1a9dbd761;
    assign coff[6024] = 64'h786f4ab4d4a5a798;
    assign coff[6025] = 64'h36814cde8c2f44ed;
    assign coff[6026] = 64'hd4a5a7988790b54c;
    assign coff[6027] = 64'h8c2f44edc97eb322;
    assign coff[6028] = 64'h73d0bb13c97eb322;
    assign coff[6029] = 64'h2b5a58688790b54c;
    assign coff[6030] = 64'hc97eb3228c2f44ed;
    assign coff[6031] = 64'h8790b54cd4a5a798;
    assign coff[6032] = 64'h6da9b28abdfc0505;
    assign coff[6033] = 64'h1edd02d683c6ceb5;
    assign coff[6034] = 64'hbdfc050592564d76;
    assign coff[6035] = 64'h83c6ceb5e122fd2a;
    assign coff[6036] = 64'h7c39314be122fd2a;
    assign coff[6037] = 64'h4203fafb92564d76;
    assign coff[6038] = 64'he122fd2a83c6ceb5;
    assign coff[6039] = 64'h92564d76bdfc0505;
    assign coff[6040] = 64'h7e940e94ecf9cafb;
    assign coff[6041] = 64'h4c0d5f37990b1d79;
    assign coff[6042] = 64'hecf9cafb816bf16c;
    assign coff[6043] = 64'h990b1d79b3f2a0c9;
    assign coff[6044] = 64'h66f4e287b3f2a0c9;
    assign coff[6045] = 64'h13063505816bf16c;
    assign coff[6046] = 64'hb3f2a0c9990b1d79;
    assign coff[6047] = 64'h816bf16cecf9cafb;
    assign coff[6048] = 64'h66aa06f3b38db1b0;
    assign coff[6049] = 64'h1289e7528159811e;
    assign coff[6050] = 64'hb38db1b09955f90d;
    assign coff[6051] = 64'h8159811eed7618ae;
    assign coff[6052] = 64'h7ea67ee2ed7618ae;
    assign coff[6053] = 64'h4c724e509955f90d;
    assign coff[6054] = 64'hed7618ae8159811e;
    assign coff[6055] = 64'h9955f90db38db1b0;
    assign coff[6056] = 64'h7c1aa8a6e0a9175e;
    assign coff[6057] = 64'h419831f39215b2d5;
    assign coff[6058] = 64'he0a9175e83e5575a;
    assign coff[6059] = 64'h9215b2d5be67ce0d;
    assign coff[6060] = 64'h6dea4d2bbe67ce0d;
    assign coff[6061] = 64'h1f56e8a283e5575a;
    assign coff[6062] = 64'hbe67ce0d9215b2d5;
    assign coff[6063] = 64'h83e5575ae0a9175e;
    assign coff[6064] = 64'h739b00adc90d19e6;
    assign coff[6065] = 64'h2ae4070a87665f96;
    assign coff[6066] = 64'hc90d19e68c64ff53;
    assign coff[6067] = 64'h87665f96d51bf8f6;
    assign coff[6068] = 64'h7899a06ad51bf8f6;
    assign coff[6069] = 64'h36f2e61a8c64ff53;
    assign coff[6070] = 64'hd51bf8f687665f96;
    assign coff[6071] = 64'h8c64ff53c90d19e6;
    assign coff[6072] = 64'h7fd562e7f97965b4;
    assign coff[6073] = 64'h55c70c4fa0fe5ce6;
    assign coff[6074] = 64'hf97965b4802a9d19;
    assign coff[6075] = 64'ha0fe5ce6aa38f3b1;
    assign coff[6076] = 64'h5f01a31aaa38f3b1;
    assign coff[6077] = 64'h06869a4c802a9d19;
    assign coff[6078] = 64'haa38f3b1a0fe5ce6;
    assign coff[6079] = 64'h802a9d19f97965b4;
    assign coff[6080] = 64'h62ca1992ae9bab60;
    assign coff[6081] = 64'h0c4d4a5d8097b030;
    assign coff[6082] = 64'hae9bab609d35e66e;
    assign coff[6083] = 64'h8097b030f3b2b5a3;
    assign coff[6084] = 64'h7f684fd0f3b2b5a3;
    assign coff[6085] = 64'h516454a09d35e66e;
    assign coff[6086] = 64'hf3b2b5a38097b030;
    assign coff[6087] = 64'h9d35e66eae9bab60;
    assign coff[6088] = 64'h7a6ab963da9bd7c7;
    assign coff[6089] = 64'h3c1f49838effa370;
    assign coff[6090] = 64'hda9bd7c78595469d;
    assign coff[6091] = 64'h8effa370c3e0b67d;
    assign coff[6092] = 64'h71005c90c3e0b67d;
    assign coff[6093] = 64'h256428398595469d;
    assign coff[6094] = 64'hc3e0b67d8effa370;
    assign coff[6095] = 64'h8595469dda9bd7c7;
    assign coff[6096] = 64'h70c51fc8c371e32d;
    assign coff[6097] = 64'h24ebe78f8570cc30;
    assign coff[6098] = 64'hc371e32d8f3ae038;
    assign coff[6099] = 64'h8570cc30db141871;
    assign coff[6100] = 64'h7a8f33d0db141871;
    assign coff[6101] = 64'h3c8e1cd38f3ae038;
    assign coff[6102] = 64'hdb1418718570cc30;
    assign coff[6103] = 64'h8f3ae038c371e32d;
    assign coff[6104] = 64'h7f5bfe9df335a6a7;
    assign coff[6105] = 64'h510330f79ce62e11;
    assign coff[6106] = 64'hf335a6a780a40163;
    assign coff[6107] = 64'h9ce62e11aefccf09;
    assign coff[6108] = 64'h6319d1efaefccf09;
    assign coff[6109] = 64'h0cca595980a40163;
    assign coff[6110] = 64'haefccf099ce62e11;
    assign coff[6111] = 64'h80a40163f335a6a7;
    assign coff[6112] = 64'h6a4aa381b8aedd86;
    assign coff[6113] = 64'h18bb155a82696ddc;
    assign coff[6114] = 64'hb8aedd8695b55c7f;
    assign coff[6115] = 64'h82696ddce744eaa6;
    assign coff[6116] = 64'h7d969224e744eaa6;
    assign coff[6117] = 64'h4751227a95b55c7f;
    assign coff[6118] = 64'he744eaa682696ddc;
    assign coff[6119] = 64'h95b55c7fb8aedd86;
    assign coff[6120] = 64'h7d7e0e1ce6c9aae5;
    assign coff[6121] = 64'h46e8a631956f8bdd;
    assign coff[6122] = 64'he6c9aae58281f1e4;
    assign coff[6123] = 64'h956f8bddb91759cf;
    assign coff[6124] = 64'h6a907423b91759cf;
    assign coff[6125] = 64'h1936551b8281f1e4;
    assign coff[6126] = 64'hb91759cf956f8bdd;
    assign coff[6127] = 64'h8281f1e4e6c9aae5;
    assign coff[6128] = 64'h7629958cceca340c;
    assign coff[6129] = 64'h30c1b2da89a65391;
    assign coff[6130] = 64'hceca340c89d66a74;
    assign coff[6131] = 64'h89a65391cf3e4d26;
    assign coff[6132] = 64'h7659ac6fcf3e4d26;
    assign coff[6133] = 64'h3135cbf489d66a74;
    assign coff[6134] = 64'hcf3e4d2689a65391;
    assign coff[6135] = 64'h89d66a74ceca340c;
    assign coff[6136] = 64'h7ffff094ffc12b0e;
    assign coff[6137] = 64'h5a5600eca5512388;
    assign coff[6138] = 64'hffc12b0e80000f6c;
    assign coff[6139] = 64'ha5512388a5a9ff14;
    assign coff[6140] = 64'h5aaedc78a5a9ff14;
    assign coff[6141] = 64'h003ed4f280000f6c;
    assign coff[6142] = 64'ha5a9ff14a5512388;
    assign coff[6143] = 64'h80000f6cffc12b0e;
    assign coff[6144] = 64'h5ac09781a5bbcf0b;
    assign coff[6145] = 64'h0057f6e980001e3a;
    assign coff[6146] = 64'ha5bbcf0ba53f687f;
    assign coff[6147] = 64'h80001e3affa80917;
    assign coff[6148] = 64'h7fffe1c6ffa80917;
    assign coff[6149] = 64'h5a4430f5a53f687f;
    assign coff[6150] = 64'hffa8091780001e3a;
    assign coff[6151] = 64'ha53f687fa5bbcf0b;
    assign coff[6152] = 64'h76633cedcf558b06;
    assign coff[6153] = 64'h314cfe7f89e0164d;
    assign coff[6154] = 64'hcf558b06899cc313;
    assign coff[6155] = 64'h89e0164dceb30181;
    assign coff[6156] = 64'h761fe9b3ceb30181;
    assign coff[6157] = 64'h30aa74fa899cc313;
    assign coff[6158] = 64'hceb3018189e0164d;
    assign coff[6159] = 64'h899cc313cf558b06;
    assign coff[6160] = 64'h6a9e5e58b92c47ae;
    assign coff[6161] = 64'h194ef88e8286e79e;
    assign coff[6162] = 64'hb92c47ae9561a1a8;
    assign coff[6163] = 64'h8286e79ee6b10772;
    assign coff[6164] = 64'h7d791862e6b10772;
    assign coff[6165] = 64'h46d3b8529561a1a8;
    assign coff[6166] = 64'he6b107728286e79e;
    assign coff[6167] = 64'h9561a1a8b92c47ae;
    assign coff[6168] = 64'h7d9b6ad3e75d93e0;
    assign coff[6169] = 64'h4765ffe695c35f53;
    assign coff[6170] = 64'he75d93e08264952d;
    assign coff[6171] = 64'h95c35f53b89a001a;
    assign coff[6172] = 64'h6a3ca0adb89a001a;
    assign coff[6173] = 64'h18a26c208264952d;
    assign coff[6174] = 64'hb89a001a95c35f53;
    assign coff[6175] = 64'h8264952de75d93e0;
    assign coff[6176] = 64'h6329b827af1045f3;
    assign coff[6177] = 64'h0ce35ae180a686c2;
    assign coff[6178] = 64'haf1045f39cd647d9;
    assign coff[6179] = 64'h80a686c2f31ca51f;
    assign coff[6180] = 64'h7f59793ef31ca51f;
    assign coff[6181] = 64'h50efba0d9cd647d9;
    assign coff[6182] = 64'hf31ca51f80a686c2;
    assign coff[6183] = 64'h9cd647d9af1045f3;
    assign coff[6184] = 64'h7a967153db2c29a9;
    assign coff[6185] = 64'h3ca440188f46c639;
    assign coff[6186] = 64'hdb2c29a985698ead;
    assign coff[6187] = 64'h8f46c639c35bbfe8;
    assign coff[6188] = 64'h70b939c7c35bbfe8;
    assign coff[6189] = 64'h24d3d65785698ead;
    assign coff[6190] = 64'hc35bbfe88f46c639;
    assign coff[6191] = 64'h85698eaddb2c29a9;
    assign coff[6192] = 64'h710c2875c3f6e7b7;
    assign coff[6193] = 64'h257c30d8859ca076;
    assign coff[6194] = 64'hc3f6e7b78ef3d78b;
    assign coff[6195] = 64'h859ca076da83cf28;
    assign coff[6196] = 64'h7a635f8ada83cf28;
    assign coff[6197] = 64'h3c0918498ef3d78b;
    assign coff[6198] = 64'hda83cf28859ca076;
    assign coff[6199] = 64'h8ef3d78bc3f6e7b7;
    assign coff[6200] = 64'h7f6ab7b8f3cbba12;
    assign coff[6201] = 64'h5177b8c29d45e389;
    assign coff[6202] = 64'hf3cbba1280954848;
    assign coff[6203] = 64'h9d45e389ae88473e;
    assign coff[6204] = 64'h62ba1c77ae88473e;
    assign coff[6205] = 64'h0c3445ee80954848;
    assign coff[6206] = 64'hae88473e9d45e389;
    assign coff[6207] = 64'h80954848f3cbba12;
    assign coff[6208] = 64'h5f1278ebaa4b9ce3;
    assign coff[6209] = 64'h069fb3c9802be796;
    assign coff[6210] = 64'haa4b9ce3a0ed8715;
    assign coff[6211] = 64'h802be796f9604c37;
    assign coff[6212] = 64'h7fd4186af9604c37;
    assign coff[6213] = 64'h55b4631da0ed8715;
    assign coff[6214] = 64'hf9604c37802be796;
    assign coff[6215] = 64'ha0ed8715aa4b9ce3;
    assign coff[6216] = 64'h78a20a03d533a7cf;
    assign coff[6217] = 64'h370998028c6fcb95;
    assign coff[6218] = 64'hd533a7cf875df5fd;
    assign coff[6219] = 64'h8c6fcb95c8f667fe;
    assign coff[6220] = 64'h7390346bc8f667fe;
    assign coff[6221] = 64'h2acc5831875df5fd;
    assign coff[6222] = 64'hc8f667fe8c6fcb95;
    assign coff[6223] = 64'h875df5fdd533a7cf;
    assign coff[6224] = 64'h6df72c30be7d6442;
    assign coff[6225] = 64'h1f6f462f83eb810a;
    assign coff[6226] = 64'hbe7d64429208d3d0;
    assign coff[6227] = 64'h83eb810ae090b9d1;
    assign coff[6228] = 64'h7c147ef6e090b9d1;
    assign coff[6229] = 64'h41829bbe9208d3d0;
    assign coff[6230] = 64'he090b9d183eb810a;
    assign coff[6231] = 64'h9208d3d0be7d6442;
    assign coff[6232] = 64'h7eaa204ced8ef72e;
    assign coff[6233] = 64'h4c86754e9964fda7;
    assign coff[6234] = 64'hed8ef72e8155dfb4;
    assign coff[6235] = 64'h9964fda7b3798ab2;
    assign coff[6236] = 64'h669b0259b3798ab2;
    assign coff[6237] = 64'h127108d28155dfb4;
    assign coff[6238] = 64'hb3798ab29964fda7;
    assign coff[6239] = 64'h8155dfb4ed8ef72e;
    assign coff[6240] = 64'h6703cf58b406d969;
    assign coff[6241] = 64'h131f0f2c816fb020;
    assign coff[6242] = 64'hb406d96998fc30a8;
    assign coff[6243] = 64'h816fb020ece0f0d4;
    assign coff[6244] = 64'h7e904fe0ece0f0d4;
    assign coff[6245] = 64'h4bf9269798fc30a8;
    assign coff[6246] = 64'hece0f0d4816fb020;
    assign coff[6247] = 64'h98fc30a8b406d969;
    assign coff[6248] = 64'h7c3f3e42e13b61e9;
    assign coff[6249] = 64'h421981f7926345e1;
    assign coff[6250] = 64'he13b61e983c0c1be;
    assign coff[6251] = 64'h926345e1bde67e09;
    assign coff[6252] = 64'h6d9cba1fbde67e09;
    assign coff[6253] = 64'h1ec49e1783c0c1be;
    assign coff[6254] = 64'hbde67e09926345e1;
    assign coff[6255] = 64'h83c0c1bee13b61e9;
    assign coff[6256] = 64'h73db6c91c99571b3;
    assign coff[6257] = 64'h2b71fd4887993ac6;
    assign coff[6258] = 64'hc99571b38c24936f;
    assign coff[6259] = 64'h87993ac6d48e02b8;
    assign coff[6260] = 64'h7866c53ad48e02b8;
    assign coff[6261] = 64'h366a8e4d8c24936f;
    assign coff[6262] = 64'hd48e02b887993ac6;
    assign coff[6263] = 64'h8c24936fc99571b3;
    assign coff[6264] = 64'h7fdcba51fa1003c8;
    assign coff[6265] = 64'h5636bdefa163aca2;
    assign coff[6266] = 64'hfa1003c8802345af;
    assign coff[6267] = 64'ha163aca2a9c94211;
    assign coff[6268] = 64'h5e9c535ea9c94211;
    assign coff[6269] = 64'h05effc38802345af;
    assign coff[6270] = 64'ha9c94211a163aca2;
    assign coff[6271] = 64'h802345affa1003c8;
    assign coff[6272] = 64'h5cf0b2afa7fcecc4;
    assign coff[6273] = 64'h037c1a22800c255a;
    assign coff[6274] = 64'ha7fcecc4a30f4d51;
    assign coff[6275] = 64'h800c255afc83e5de;
    assign coff[6276] = 64'h7ff3daa6fc83e5de;
    assign coff[6277] = 64'h5803133ca30f4d51;
    assign coff[6278] = 64'hfc83e5de800c255a;
    assign coff[6279] = 64'ha30f4d51a7fcecc4;
    assign coff[6280] = 64'h778bdb19d241127a;
    assign coff[6281] = 64'h342f51498b1eedf4;
    assign coff[6282] = 64'hd241127a887424e7;
    assign coff[6283] = 64'h8b1eedf4cbd0aeb7;
    assign coff[6284] = 64'h74e1120ccbd0aeb7;
    assign coff[6285] = 64'h2dbeed86887424e7;
    assign coff[6286] = 64'hcbd0aeb78b1eedf4;
    assign coff[6287] = 64'h887424e7d241127a;
    assign coff[6288] = 64'h6c531f67bbcf940a;
    assign coff[6289] = 64'h1c614f8b832f94b8;
    assign coff[6290] = 64'hbbcf940a93ace099;
    assign coff[6291] = 64'h832f94b8e39eb075;
    assign coff[6292] = 64'h7cd06b48e39eb075;
    assign coff[6293] = 64'h44306bf693ace099;
    assign coff[6294] = 64'he39eb075832f94b8;
    assign coff[6295] = 64'h93ace099bbcf940a;
    assign coff[6296] = 64'h7e2c8002ea749c47;
    assign coff[6297] = 64'h49fbeeea978c20c8;
    assign coff[6298] = 64'hea749c4781d37ffe;
    assign coff[6299] = 64'h978c20c8b6041116;
    assign coff[6300] = 64'h6873df38b6041116;
    assign coff[6301] = 64'h158b63b981d37ffe;
    assign coff[6302] = 64'hb6041116978c20c8;
    assign coff[6303] = 64'h81d37ffeea749c47;
    assign coff[6304] = 64'h651e8faab18582a8;
    assign coff[6305] = 64'h10027107810150ca;
    assign coff[6306] = 64'hb18582a89ae17056;
    assign coff[6307] = 64'h810150caeffd8ef9;
    assign coff[6308] = 64'h7efeaf36effd8ef9;
    assign coff[6309] = 64'h4e7a7d589ae17056;
    assign coff[6310] = 64'heffd8ef9810150ca;
    assign coff[6311] = 64'h9ae17056b18582a8;
    assign coff[6312] = 64'h7b745c91de312a7a;
    assign coff[6313] = 64'h3f63c43b90cc7322;
    assign coff[6314] = 64'hde312a7a848ba36f;
    assign coff[6315] = 64'h90cc7322c09c3bc5;
    assign coff[6316] = 64'h6f338cdec09c3bc5;
    assign coff[6317] = 64'h21ced586848ba36f;
    assign coff[6318] = 64'hc09c3bc590cc7322;
    assign coff[6319] = 64'h848ba36fde312a7a;
    assign coff[6320] = 64'h727c9e47c6c1c2d4;
    assign coff[6321] = 64'h287a3604869190c7;
    assign coff[6322] = 64'hc6c1c2d48d8361b9;
    assign coff[6323] = 64'h869190c7d785c9fc;
    assign coff[6324] = 64'h796e6f39d785c9fc;
    assign coff[6325] = 64'h393e3d2c8d8361b9;
    assign coff[6326] = 64'hd785c9fc869190c7;
    assign coff[6327] = 64'h8d8361b9c6c1c2d4;
    assign coff[6328] = 64'h7fad9127f6ed2bd4;
    assign coff[6329] = 64'h53ddb2b69f4d5371;
    assign coff[6330] = 64'hf6ed2bd480526ed9;
    assign coff[6331] = 64'h9f4d5371ac224d4a;
    assign coff[6332] = 64'h60b2ac8fac224d4a;
    assign coff[6333] = 64'h0912d42c80526ed9;
    assign coff[6334] = 64'hac224d4a9f4d5371;
    assign coff[6335] = 64'h80526ed9f6ed2bd4;
    assign coff[6336] = 64'h6125960aaca78453;
    assign coff[6337] = 64'h09c247f5805f6009;
    assign coff[6338] = 64'haca784539eda69f6;
    assign coff[6339] = 64'h805f6009f63db80b;
    assign coff[6340] = 64'h7fa09ff7f63db80b;
    assign coff[6341] = 64'h53587bad9eda69f6;
    assign coff[6342] = 64'hf63db80b805f6009;
    assign coff[6343] = 64'h9eda69f6aca78453;
    assign coff[6344] = 64'h79a59ec3d82cd6aa;
    assign coff[6345] = 64'h39db620b8dd27b3c;
    assign coff[6346] = 64'hd82cd6aa865a613d;
    assign coff[6347] = 64'h8dd27b3cc6249df5;
    assign coff[6348] = 64'h722d84c4c6249df5;
    assign coff[6349] = 64'h27d32956865a613d;
    assign coff[6350] = 64'hc6249df58dd27b3c;
    assign coff[6351] = 64'h865a613dd82cd6aa;
    assign coff[6352] = 64'h6f8a43edc1354e97;
    assign coff[6353] = 64'h227863e584ba8f98;
    assign coff[6354] = 64'hc1354e979075bc13;
    assign coff[6355] = 64'h84ba8f98dd879c1b;
    assign coff[6356] = 64'h7b457068dd879c1b;
    assign coff[6357] = 64'h3ecab1699075bc13;
    assign coff[6358] = 64'hdd879c1b84ba8f98;
    assign coff[6359] = 64'h9075bc13c1354e97;
    assign coff[6360] = 64'h7f143852f0ac2a16;
    assign coff[6361] = 64'h4f052ec09b4dad06;
    assign coff[6362] = 64'hf0ac2a1680ebc7ae;
    assign coff[6363] = 64'h9b4dad06b0fad140;
    assign coff[6364] = 64'h64b252fab0fad140;
    assign coff[6365] = 64'h0f53d5ea80ebc7ae;
    assign coff[6366] = 64'hb0fad1409b4dad06;
    assign coff[6367] = 64'h80ebc7aef0ac2a16;
    assign coff[6368] = 64'h68d92c5db693e752;
    assign coff[6369] = 64'h1638ba7a81f193be;
    assign coff[6370] = 64'hb693e7529726d3a3;
    assign coff[6371] = 64'h81f193bee9c74586;
    assign coff[6372] = 64'h7e0e6c42e9c74586;
    assign coff[6373] = 64'h496c18ae9726d3a3;
    assign coff[6374] = 64'he9c7458681f193be;
    assign coff[6375] = 64'h9726d3a3b693e752;
    assign coff[6376] = 64'h7cf6f720e44a57f4;
    assign coff[6377] = 64'h44c50e53940affb9;
    assign coff[6378] = 64'he44a57f4830908e0;
    assign coff[6379] = 64'h940affb9bb3af1ad;
    assign coff[6380] = 64'h6bf50047bb3af1ad;
    assign coff[6381] = 64'h1bb5a80c830908e0;
    assign coff[6382] = 64'hbb3af1ad940affb9;
    assign coff[6383] = 64'h830908e0e44a57f4;
    assign coff[6384] = 64'h75285d3bcc7184ba;
    assign coff[6385] = 64'h2e63117c88b375ca;
    assign coff[6386] = 64'hcc7184ba8ad7a2c5;
    assign coff[6387] = 64'h88b375cad19cee84;
    assign coff[6388] = 64'h774c8a36d19cee84;
    assign coff[6389] = 64'h338e7b468ad7a2c5;
    assign coff[6390] = 64'hd19cee8488b375ca;
    assign coff[6391] = 64'h8ad7a2c5cc7184ba;
    assign coff[6392] = 64'h7ff82beffd33c61f;
    assign coff[6393] = 64'h58827dbea3889cb8;
    assign coff[6394] = 64'hfd33c61f8007d411;
    assign coff[6395] = 64'ha3889cb8a77d8242;
    assign coff[6396] = 64'h5c776348a77d8242;
    assign coff[6397] = 64'h02cc39e18007d411;
    assign coff[6398] = 64'ha77d8242a3889cb8;
    assign coff[6399] = 64'h8007d411fd33c61f;
    assign coff[6400] = 64'h5bda6a5da6daa5fe;
    assign coff[6401] = 64'h01ea11f78003aa36;
    assign coff[6402] = 64'ha6daa5fea42595a3;
    assign coff[6403] = 64'h8003aa36fe15ee09;
    assign coff[6404] = 64'h7ffc55cafe15ee09;
    assign coff[6405] = 64'h59255a02a42595a3;
    assign coff[6406] = 64'hfe15ee098003aa36;
    assign coff[6407] = 64'ha42595a3a6daa5fe;
    assign coff[6408] = 64'h76f9d721d0ca65c9;
    assign coff[6409] = 64'h32bf22508a7d3e3e;
    assign coff[6410] = 64'hd0ca65c9890628df;
    assign coff[6411] = 64'h8a7d3e3ecd40ddb0;
    assign coff[6412] = 64'h7582c1c2cd40ddb0;
    assign coff[6413] = 64'h2f359a37890628df;
    assign coff[6414] = 64'hcd40ddb08a7d3e3e;
    assign coff[6415] = 64'h890628dfd0ca65c9;
    assign coff[6416] = 64'h6b7ad142ba7c96d4;
    assign coff[6417] = 64'h1ad8a88782d8d492;
    assign coff[6418] = 64'hba7c96d494852ebe;
    assign coff[6419] = 64'h82d8d492e5275779;
    assign coff[6420] = 64'h7d272b6ee5275779;
    assign coff[6421] = 64'h4583692c94852ebe;
    assign coff[6422] = 64'he527577982d8d492;
    assign coff[6423] = 64'h94852ebeba7c96d4;
    assign coff[6424] = 64'h7de662b3e8e8a621;
    assign coff[6425] = 64'h48b25e2596a5b82a;
    assign coff[6426] = 64'he8e8a62182199d4d;
    assign coff[6427] = 64'h96a5b82ab74da1db;
    assign coff[6428] = 64'h695a47d6b74da1db;
    assign coff[6429] = 64'h171759df82199d4d;
    assign coff[6430] = 64'hb74da1db96a5b82a;
    assign coff[6431] = 64'h82199d4de8e8a621;
    assign coff[6432] = 64'h6426121eb0495af0;
    assign coff[6433] = 64'h0e732d4280d1782a;
    assign coff[6434] = 64'hb0495af09bd9ede2;
    assign coff[6435] = 64'h80d1782af18cd2be;
    assign coff[6436] = 64'h7f2e87d6f18cd2be;
    assign coff[6437] = 64'h4fb6a5109bd9ede2;
    assign coff[6438] = 64'hf18cd2be80d1782a;
    assign coff[6439] = 64'h9bd9ede2b0495af0;
    assign coff[6440] = 64'h7b07c612dcadfbc5;
    assign coff[6441] = 64'h3e05343790077422;
    assign coff[6442] = 64'hdcadfbc584f839ee;
    assign coff[6443] = 64'h90077422c1facbc9;
    assign coff[6444] = 64'h6ff88bdec1facbc9;
    assign coff[6445] = 64'h2352043b84f839ee;
    assign coff[6446] = 64'hc1facbc990077422;
    assign coff[6447] = 64'h84f839eedcadfbc5;
    assign coff[6448] = 64'h71c694d2c55b33e2;
    assign coff[6449] = 64'h26fbf3ce8614befb;
    assign coff[6450] = 64'hc55b33e28e396b2e;
    assign coff[6451] = 64'h8614befbd9040c32;
    assign coff[6452] = 64'h79eb4105d9040c32;
    assign coff[6453] = 64'h3aa4cc1e8e396b2e;
    assign coff[6454] = 64'hd9040c328614befb;
    assign coff[6455] = 64'h8e396b2ec55b33e2;
    assign coff[6456] = 64'h7f8e99e6f55c3e72;
    assign coff[6457] = 64'h52ac4db49e47b944;
    assign coff[6458] = 64'hf55c3e728071661a;
    assign coff[6459] = 64'h9e47b944ad53b24c;
    assign coff[6460] = 64'h61b846bcad53b24c;
    assign coff[6461] = 64'h0aa3c18e8071661a;
    assign coff[6462] = 64'had53b24c9e47b944;
    assign coff[6463] = 64'h8071661af55c3e72;
    assign coff[6464] = 64'h601de1caab77ef77;
    assign coff[6465] = 64'h0831264c80432d75;
    assign coff[6466] = 64'hab77ef779fe21e36;
    assign coff[6467] = 64'h80432d75f7ced9b4;
    assign coff[6468] = 64'h7fbcd28bf7ced9b4;
    assign coff[6469] = 64'h548810899fe21e36;
    assign coff[6470] = 64'hf7ced9b480432d75;
    assign coff[6471] = 64'h9fe21e36ab77ef77;
    assign coff[6472] = 64'h79262a3ad6af735c;
    assign coff[6473] = 64'h387393998d1eec83;
    assign coff[6474] = 64'hd6af735c86d9d5c6;
    assign coff[6475] = 64'h8d1eec83c78c6c67;
    assign coff[6476] = 64'h72e1137dc78c6c67;
    assign coff[6477] = 64'h29508ca486d9d5c6;
    assign coff[6478] = 64'hc78c6c678d1eec83;
    assign coff[6479] = 64'h86d9d5c6d6af735c;
    assign coff[6480] = 64'h6ec2daa2bfd81cd5;
    assign coff[6481] = 64'h20f477aa8450a5f7;
    assign coff[6482] = 64'hbfd81cd5913d255e;
    assign coff[6483] = 64'h8450a5f7df0b8856;
    assign coff[6484] = 64'h7baf5a09df0b8856;
    assign coff[6485] = 64'h4027e32b913d255e;
    assign coff[6486] = 64'hdf0b88568450a5f7;
    assign coff[6487] = 64'h913d255ebfd81cd5;
    assign coff[6488] = 64'h7ee19e6fef1d3d4e;
    assign coff[6489] = 64'h4dc751d89a575fae;
    assign coff[6490] = 64'hef1d3d4e811e6191;
    assign coff[6491] = 64'h9a575faeb238ae28;
    assign coff[6492] = 64'h65a8a052b238ae28;
    assign coff[6493] = 64'h10e2c2b2811e6191;
    assign coff[6494] = 64'hb238ae289a575fae;
    assign coff[6495] = 64'h811e6191ef1d3d4e;
    assign coff[6496] = 64'h67f07ec5b54befba;
    assign coff[6497] = 64'h14ac4ad781ae3294;
    assign coff[6498] = 64'hb54befba980f813b;
    assign coff[6499] = 64'h81ae3294eb53b529;
    assign coff[6500] = 64'h7e51cd6ceb53b529;
    assign coff[6501] = 64'h4ab41046980f813b;
    assign coff[6502] = 64'heb53b52981ae3294;
    assign coff[6503] = 64'h980f813bb54befba;
    assign coff[6504] = 64'h7c9d81a3e2c24ca2;
    assign coff[6505] = 64'h437094f1933509f0;
    assign coff[6506] = 64'he2c24ca283627e5d;
    assign coff[6507] = 64'h933509f0bc8f6b0f;
    assign coff[6508] = 64'h6ccaf610bc8f6b0f;
    assign coff[6509] = 64'h1d3db35e83627e5d;
    assign coff[6510] = 64'hbc8f6b0f933509f0;
    assign coff[6511] = 64'h83627e5de2c24ca2;
    assign coff[6512] = 64'h748423e0cb0275b8;
    assign coff[6513] = 64'h2ceb650d882408ce;
    assign coff[6514] = 64'hcb0275b88b7bdc20;
    assign coff[6515] = 64'h882408ced3149af3;
    assign coff[6516] = 64'h77dbf732d3149af3;
    assign coff[6517] = 64'h34fd8a488b7bdc20;
    assign coff[6518] = 64'hd3149af3882408ce;
    assign coff[6519] = 64'h8b7bdc20cb0275b8;
    assign coff[6520] = 64'h7fecea67fba1cf66;
    assign coff[6521] = 64'h575e4cfaa274570d;
    assign coff[6522] = 64'hfba1cf6680131599;
    assign coff[6523] = 64'ha274570da8a1b306;
    assign coff[6524] = 64'h5d8ba8f3a8a1b306;
    assign coff[6525] = 64'h045e309a80131599;
    assign coff[6526] = 64'ha8a1b306a274570d;
    assign coff[6527] = 64'h80131599fba1cf66;
    assign coff[6528] = 64'h5e0365bba922982c;
    assign coff[6529] = 64'h050dffe780198f50;
    assign coff[6530] = 64'ha922982ca1fc9a45;
    assign coff[6531] = 64'h80198f50faf20019;
    assign coff[6532] = 64'h7fe670b0faf20019;
    assign coff[6533] = 64'h56dd67d4a1fc9a45;
    assign coff[6534] = 64'hfaf2001980198f50;
    assign coff[6535] = 64'ha1fc9a45a922982c;
    assign coff[6536] = 64'h78194336d3b982a8;
    assign coff[6537] = 64'h359d7d398bc51f34;
    assign coff[6538] = 64'hd3b982a887e6bcca;
    assign coff[6539] = 64'h8bc51f34ca6282c7;
    assign coff[6540] = 64'h743ae0ccca6282c7;
    assign coff[6541] = 64'h2c467d5887e6bcca;
    assign coff[6542] = 64'hca6282c78bc51f34;
    assign coff[6543] = 64'h87e6bccad3b982a8;
    assign coff[6544] = 64'h6d274070bd25323d;
    assign coff[6545] = 64'h1de8de75838b24b8;
    assign coff[6546] = 64'hbd25323d92d8bf90;
    assign coff[6547] = 64'h838b24b8e217218b;
    assign coff[6548] = 64'h7c74db48e217218b;
    assign coff[6549] = 64'h42dacdc392d8bf90;
    assign coff[6550] = 64'he217218b838b24b8;
    assign coff[6551] = 64'h92d8bf90bd25323d;
    assign coff[6552] = 64'h7e6dc00cec01670f;
    assign coff[6553] = 64'h4b42a5809876904a;
    assign coff[6554] = 64'hec01670f81923ff4;
    assign coff[6555] = 64'h9876904ab4bd5a80;
    assign coff[6556] = 64'h67896fb6b4bd5a80;
    assign coff[6557] = 64'h13fe98f181923ff4;
    assign coff[6558] = 64'hb4bd5a809876904a;
    assign coff[6559] = 64'h81923ff4ec01670f;
    assign coff[6560] = 64'h66132738b2c4b0ea;
    assign coff[6561] = 64'h119116c981360ec9;
    assign coff[6562] = 64'hb2c4b0ea99ecd8c8;
    assign coff[6563] = 64'h81360ec9ee6ee937;
    assign coff[6564] = 64'h7ec9f137ee6ee937;
    assign coff[6565] = 64'h4d3b4f1699ecd8c8;
    assign coff[6566] = 64'hee6ee93781360ec9;
    assign coff[6567] = 64'h99ecd8c8b2c4b0ea;
    assign coff[6568] = 64'h7bdc30a1dfb5a6d9;
    assign coff[6569] = 64'h40bfe29f9195bba3;
    assign coff[6570] = 64'hdfb5a6d98423cf5f;
    assign coff[6571] = 64'h9195bba3bf401d61;
    assign coff[6572] = 64'h6e6a445dbf401d61;
    assign coff[6573] = 64'h204a59278423cf5f;
    assign coff[6574] = 64'hbf401d619195bba3;
    assign coff[6575] = 64'h8423cf5fdfb5a6d9;
    assign coff[6576] = 64'h732e3dcfc82a86bd;
    assign coff[6577] = 64'h29f6e8bb8713110a;
    assign coff[6578] = 64'hc82a86bd8cd1c231;
    assign coff[6579] = 64'h8713110ad6091745;
    assign coff[6580] = 64'h78eceef6d6091745;
    assign coff[6581] = 64'h37d579438cd1c231;
    assign coff[6582] = 64'hd60917458713110a;
    assign coff[6583] = 64'h8cd1c231c82a86bd;
    assign coff[6584] = 64'h7fc79c4bf87e72c4;
    assign coff[6585] = 64'h550bdc01a056a7f9;
    assign coff[6586] = 64'hf87e72c4803863b5;
    assign coff[6587] = 64'ha056a7f9aaf423ff;
    assign coff[6588] = 64'h5fa95807aaf423ff;
    assign coff[6589] = 64'h07818d3c803863b5;
    assign coff[6590] = 64'haaf423ffa056a7f9;
    assign coff[6591] = 64'h803863b5f87e72c4;
    assign coff[6592] = 64'h62298b81adda4fc3;
    assign coff[6593] = 64'h0b53094d80807e3a;
    assign coff[6594] = 64'hadda4fc39dd6747f;
    assign coff[6595] = 64'h80807e3af4acf6b3;
    assign coff[6596] = 64'h7f7f81c6f4acf6b3;
    assign coff[6597] = 64'h5225b03d9dd6747f;
    assign coff[6598] = 64'hf4acf6b380807e3a;
    assign coff[6599] = 64'h9dd6747fadda4fc3;
    assign coff[6600] = 64'h7a2062b5d9abc305;
    assign coff[6601] = 64'h3b40f5798e8a70d7;
    assign coff[6602] = 64'hd9abc30585df9d4b;
    assign coff[6603] = 64'h8e8a70d7c4bf0a87;
    assign coff[6604] = 64'h71758f29c4bf0a87;
    assign coff[6605] = 64'h26543cfb85df9d4b;
    assign coff[6606] = 64'hc4bf0a878e8a70d7;
    assign coff[6607] = 64'h85df9d4bd9abc305;
    assign coff[6608] = 64'h704d6060c294ec12;
    assign coff[6609] = 64'h23fafbec852939da;
    assign coff[6610] = 64'hc294ec128fb29fa0;
    assign coff[6611] = 64'h852939dadc050414;
    assign coff[6612] = 64'h7ad6c626dc050414;
    assign coff[6613] = 64'h3d6b13ee8fb29fa0;
    assign coff[6614] = 64'hdc050414852939da;
    assign coff[6615] = 64'h8fb29fa0c294ec12;
    assign coff[6616] = 64'h7f41ec01f23bae24;
    assign coff[6617] = 64'h503fffc49c47dc31;
    assign coff[6618] = 64'hf23bae2480be13ff;
    assign coff[6619] = 64'h9c47dc31afc0003c;
    assign coff[6620] = 64'h63b823cfafc0003c;
    assign coff[6621] = 64'h0dc451dc80be13ff;
    assign coff[6622] = 64'hafc0003c9c47dc31;
    assign coff[6623] = 64'h80be13fff23bae24;
    assign coff[6624] = 64'h69bdcf29b7deb38f;
    assign coff[6625] = 64'h17c44ecd8239d104;
    assign coff[6626] = 64'hb7deb38f964230d7;
    assign coff[6627] = 64'h8239d104e83bb133;
    assign coff[6628] = 64'h7dc62efce83bb133;
    assign coff[6629] = 64'h48214c71964230d7;
    assign coff[6630] = 64'he83bb1338239d104;
    assign coff[6631] = 64'h964230d7b7deb38f;
    assign coff[6632] = 64'h7d4b9b46e5d374c1;
    assign coff[6633] = 64'h4616e0fc94e51efd;
    assign coff[6634] = 64'he5d374c182b464ba;
    assign coff[6635] = 64'h94e51efdb9e91f04;
    assign coff[6636] = 64'h6b1ae103b9e91f04;
    assign coff[6637] = 64'h1a2c8b3f82b464ba;
    assign coff[6638] = 64'hb9e91f0494e51efd;
    assign coff[6639] = 64'h82b464bae5d374c1;
    assign coff[6640] = 64'h75c8124dcde29092;
    assign coff[6641] = 64'h2fd8f41b89477c30;
    assign coff[6642] = 64'hcde290928a37edb3;
    assign coff[6643] = 64'h89477c30d0270be5;
    assign coff[6644] = 64'h76b883d0d0270be5;
    assign coff[6645] = 64'h321d6f6e8a37edb3;
    assign coff[6646] = 64'hd0270be589477c30;
    assign coff[6647] = 64'h8a37edb3cde29092;
    assign coff[6648] = 64'h7ffe7e79fec5d876;
    assign coff[6649] = 64'h59a344f6a4a072fa;
    assign coff[6650] = 64'hfec5d87680018187;
    assign coff[6651] = 64'ha4a072faa65cbb0a;
    assign coff[6652] = 64'h5b5f8d06a65cbb0a;
    assign coff[6653] = 64'h013a278a80018187;
    assign coff[6654] = 64'ha65cbb0aa4a072fa;
    assign coff[6655] = 64'h80018187fec5d876;
    assign coff[6656] = 64'h5b4df193a64acbd9;
    assign coff[6657] = 64'h012105d580014650;
    assign coff[6658] = 64'ha64acbd9a4b20e6d;
    assign coff[6659] = 64'h80014650fedefa2b;
    assign coff[6660] = 64'h7ffeb9b0fedefa2b;
    assign coff[6661] = 64'h59b53427a4b20e6d;
    assign coff[6662] = 64'hfedefa2b80014650;
    assign coff[6663] = 64'ha4b20e6da64acbd9;
    assign coff[6664] = 64'h76af1c72d00fbd43;
    assign coff[6665] = 64'h32064e1e8a2e18eb;
    assign coff[6666] = 64'hd00fbd438950e38e;
    assign coff[6667] = 64'h8a2e18ebcdf9b1e2;
    assign coff[6668] = 64'h75d1e715cdf9b1e2;
    assign coff[6669] = 64'h2ff042bd8950e38e;
    assign coff[6670] = 64'hcdf9b1e28a2e18eb;
    assign coff[6671] = 64'h8950e38ed00fbd43;
    assign coff[6672] = 64'h6b0d1bdfb9d418af;
    assign coff[6673] = 64'h1a13f0b682af437e;
    assign coff[6674] = 64'hb9d418af94f2e421;
    assign coff[6675] = 64'h82af437ee5ec0f4a;
    assign coff[6676] = 64'h7d50bc82e5ec0f4a;
    assign coff[6677] = 64'h462be75194f2e421;
    assign coff[6678] = 64'he5ec0f4a82af437e;
    assign coff[6679] = 64'h94f2e421b9d418af;
    assign coff[6680] = 64'h7dc181e8e822ff90;
    assign coff[6681] = 64'h480c87e896340939;
    assign coff[6682] = 64'he822ff90823e7e18;
    assign coff[6683] = 64'h96340939b7f37818;
    assign coff[6684] = 64'h69cbf6c7b7f37818;
    assign coff[6685] = 64'h17dd0070823e7e18;
    assign coff[6686] = 64'hb7f3781896340939;
    assign coff[6687] = 64'h823e7e18e822ff90;
    assign coff[6688] = 64'h63a86015afac6d58;
    assign coff[6689] = 64'h0dab54ef80bb6274;
    assign coff[6690] = 64'hafac6d589c579feb;
    assign coff[6691] = 64'h80bb6274f254ab11;
    assign coff[6692] = 64'h7f449d8cf254ab11;
    assign coff[6693] = 64'h505392a89c579feb;
    assign coff[6694] = 64'hf254ab1180bb6274;
    assign coff[6695] = 64'h9c579febafac6d58;
    assign coff[6696] = 64'h7acfb336dbece636;
    assign coff[6697] = 64'h3d5505d28fa69293;
    assign coff[6698] = 64'hdbece63685304cca;
    assign coff[6699] = 64'h8fa69293c2aafa2e;
    assign coff[6700] = 64'h70596d6dc2aafa2e;
    assign coff[6701] = 64'h241319ca85304cca;
    assign coff[6702] = 64'hc2aafa2e8fa69293;
    assign coff[6703] = 64'h85304ccadbece636;
    assign coff[6704] = 64'h7169ea8fc4a8c497;
    assign coff[6705] = 64'h263c417f85d81905;
    assign coff[6706] = 64'hc4a8c4978e961571;
    assign coff[6707] = 64'h85d81905d9c3be81;
    assign coff[6708] = 64'h7a27e6fbd9c3be81;
    assign coff[6709] = 64'h3b573b698e961571;
    assign coff[6710] = 64'hd9c3be8185d81905;
    assign coff[6711] = 64'h8e961571c4a8c497;
    assign coff[6712] = 64'h7f7d4617f493ee2b;
    assign coff[6713] = 64'h5212687b9dc65539;
    assign coff[6714] = 64'hf493ee2b8082b9e9;
    assign coff[6715] = 64'h9dc65539aded9785;
    assign coff[6716] = 64'h6239aac7aded9785;
    assign coff[6717] = 64'h0b6c11d58082b9e9;
    assign coff[6718] = 64'haded97859dc65539;
    assign coff[6719] = 64'h8082b9e9f493ee2b;
    assign coff[6720] = 64'h5f98a34aaae15d2a;
    assign coff[6721] = 64'h0768762e8036ece0;
    assign coff[6722] = 64'haae15d2aa0675cb6;
    assign coff[6723] = 64'h8036ece0f89789d2;
    assign coff[6724] = 64'h7fc91320f89789d2;
    assign coff[6725] = 64'h551ea2d6a0675cb6;
    assign coff[6726] = 64'hf89789d28036ece0;
    assign coff[6727] = 64'ha0675cb6aae15d2a;
    assign coff[6728] = 64'h78e4af44d5f159b3;
    assign coff[6729] = 64'h37beda938cc6cde5;
    assign coff[6730] = 64'hd5f159b3871b50bc;
    assign coff[6731] = 64'h8cc6cde5c841256d;
    assign coff[6732] = 64'h7339321bc841256d;
    assign coff[6733] = 64'h2a0ea64d871b50bc;
    assign coff[6734] = 64'hc841256d8cc6cde5;
    assign coff[6735] = 64'h871b50bcd5f159b3;
    assign coff[6736] = 64'h6e5d8b91bf2a708f;
    assign coff[6737] = 64'h203206a4841d7aaa;
    assign coff[6738] = 64'hbf2a708f91a2746f;
    assign coff[6739] = 64'h841d7aaadfcdf95c;
    assign coff[6740] = 64'h7be28556dfcdf95c;
    assign coff[6741] = 64'h40d58f7191a2746f;
    assign coff[6742] = 64'hdfcdf95c841d7aaa;
    assign coff[6743] = 64'h91a2746fbf2a708f;
    assign coff[6744] = 64'h7ec67bc5ee560473;
    assign coff[6745] = 64'h4d2742c299ddb0aa;
    assign coff[6746] = 64'hee5604738139843b;
    assign coff[6747] = 64'h99ddb0aab2d8bd3e;
    assign coff[6748] = 64'h66224f56b2d8bd3e;
    assign coff[6749] = 64'h11a9fb8d8139843b;
    assign coff[6750] = 64'hb2d8bd3e99ddb0aa;
    assign coff[6751] = 64'h8139843bee560473;
    assign coff[6752] = 64'h677aa6b8b4a9079f;
    assign coff[6753] = 64'h13e5c58e818e555c;
    assign coff[6754] = 64'hb4a9079f98855948;
    assign coff[6755] = 64'h818e555cec1a3a72;
    assign coff[6756] = 64'h7e71aaa4ec1a3a72;
    assign coff[6757] = 64'h4b56f86198855948;
    assign coff[6758] = 64'hec1a3a72818e555c;
    assign coff[6759] = 64'h98855948b4a9079f;
    assign coff[6760] = 64'h7c6ef976e1feb241;
    assign coff[6761] = 64'h42c55dd492cba12f;
    assign coff[6762] = 64'he1feb2418391068a;
    assign coff[6763] = 64'h92cba12fbd3aa22c;
    assign coff[6764] = 64'h6d345ed1bd3aa22c;
    assign coff[6765] = 64'h1e014dbf8391068a;
    assign coff[6766] = 64'hbd3aa22c92cba12f;
    assign coff[6767] = 64'h8391068ae1feb241;
    assign coff[6768] = 64'h74305790ca4bb174;
    assign coff[6769] = 64'h2c2ee7ad87de0d95;
    assign coff[6770] = 64'hca4bb1748bcfa870;
    assign coff[6771] = 64'h87de0d95d3d11853;
    assign coff[6772] = 64'h7821f26bd3d11853;
    assign coff[6773] = 64'h35b44e8c8bcfa870;
    assign coff[6774] = 64'hd3d1185387de0d95;
    assign coff[6775] = 64'h8bcfa870ca4bb174;
    assign coff[6776] = 64'h7fe57025fad8e33c;
    assign coff[6777] = 64'h56caf088a1eb8dc7;
    assign coff[6778] = 64'hfad8e33c801a8fdb;
    assign coff[6779] = 64'ha1eb8dc7a9350f78;
    assign coff[6780] = 64'h5e147239a9350f78;
    assign coff[6781] = 64'h05271cc4801a8fdb;
    assign coff[6782] = 64'ha9350f78a1eb8dc7;
    assign coff[6783] = 64'h801a8fdbfad8e33c;
    assign coff[6784] = 64'h5d7a7f88a88f5698;
    assign coff[6785] = 64'h0445124980123c82;
    assign coff[6786] = 64'ha88f5698a2858078;
    assign coff[6787] = 64'h80123c82fbbaedb7;
    assign coff[6788] = 64'h7fedc37efbbaedb7;
    assign coff[6789] = 64'h5770a968a2858078;
    assign coff[6790] = 64'hfbbaedb780123c82;
    assign coff[6791] = 64'ha2858078a88f5698;
    assign coff[6792] = 64'h77d322fcd2fd1309;
    assign coff[6793] = 64'h34e6a8858b7176c8;
    assign coff[6794] = 64'hd2fd1309882cdd04;
    assign coff[6795] = 64'h8b7176c8cb19577b;
    assign coff[6796] = 64'h748e8938cb19577b;
    assign coff[6797] = 64'h2d02ecf7882cdd04;
    assign coff[6798] = 64'hcb19577b8b7176c8;
    assign coff[6799] = 64'h882cdd04d2fd1309;
    assign coff[6800] = 64'h6cbdb613bc7a0fd6;
    assign coff[6801] = 64'h1d253af5835cc2f4;
    assign coff[6802] = 64'hbc7a0fd6934249ed;
    assign coff[6803] = 64'h835cc2f4e2dac50b;
    assign coff[6804] = 64'h7ca33d0ce2dac50b;
    assign coff[6805] = 64'h4385f02a934249ed;
    assign coff[6806] = 64'he2dac50b835cc2f4;
    assign coff[6807] = 64'h934249edbc7a0fd6;
    assign coff[6808] = 64'h7e4dbbd9eb3ae80c;
    assign coff[6809] = 64'h4a9fa6459800d83c;
    assign coff[6810] = 64'heb3ae80c81b24427;
    assign coff[6811] = 64'h9800d83cb56059bb;
    assign coff[6812] = 64'h67ff27c4b56059bb;
    assign coff[6813] = 64'h14c517f481b24427;
    assign coff[6814] = 64'hb56059bb9800d83c;
    assign coff[6815] = 64'h81b24427eb3ae80c;
    assign coff[6816] = 64'h659958c9b224b9bc;
    assign coff[6817] = 64'h10c9d89e811b133d;
    assign coff[6818] = 64'hb224b9bc9a66a737;
    assign coff[6819] = 64'h811b133def362762;
    assign coff[6820] = 64'h7ee4ecc3ef362762;
    assign coff[6821] = 64'h4ddb46449a66a737;
    assign coff[6822] = 64'hef362762811b133d;
    assign coff[6823] = 64'h9a66a737b224b9bc;
    assign coff[6824] = 64'h7ba8df28def33fe3;
    assign coff[6825] = 64'h4012227891308eae;
    assign coff[6826] = 64'hdef33fe3845720d8;
    assign coff[6827] = 64'h91308eaebfeddd88;
    assign coff[6828] = 64'h6ecf7152bfeddd88;
    assign coff[6829] = 64'h210cc01d845720d8;
    assign coff[6830] = 64'hbfeddd8891308eae;
    assign coff[6831] = 64'h845720d8def33fe3;
    assign coff[6832] = 64'h72d5fbb7c775df08;
    assign coff[6833] = 64'h2938c23a86d1bb69;
    assign coff[6834] = 64'hc775df088d2a0449;
    assign coff[6835] = 64'h86d1bb69d6c73dc6;
    assign coff[6836] = 64'h792e4497d6c73dc6;
    assign coff[6837] = 64'h388a20f88d2a0449;
    assign coff[6838] = 64'hd6c73dc686d1bb69;
    assign coff[6839] = 64'h8d2a0449c775df08;
    assign coff[6840] = 64'h7fbb344ef7b5c512;
    assign coff[6841] = 64'h54752f8d9fd1870c;
    assign coff[6842] = 64'hf7b5c5128044cbb2;
    assign coff[6843] = 64'h9fd1870cab8ad073;
    assign coff[6844] = 64'h602e78f4ab8ad073;
    assign coff[6845] = 64'h084a3aee8044cbb2;
    assign coff[6846] = 64'hab8ad0739fd1870c;
    assign coff[6847] = 64'h8044cbb2f7b5c512;
    assign coff[6848] = 64'h61a80940ad4083f5;
    assign coff[6849] = 64'h0a8ab5a2806f51c1;
    assign coff[6850] = 64'had4083f59e57f6c0;
    assign coff[6851] = 64'h806f51c1f5754a5e;
    assign coff[6852] = 64'h7f90ae3ff5754a5e;
    assign coff[6853] = 64'h52bf7c0b9e57f6c0;
    assign coff[6854] = 64'hf5754a5e806f51c1;
    assign coff[6855] = 64'h9e57f6c0ad4083f5;
    assign coff[6856] = 64'h79e3971cd8ec1ca1;
    assign coff[6857] = 64'h3a8e74008e2de99e;
    assign coff[6858] = 64'hd8ec1ca1861c68e4;
    assign coff[6859] = 64'h8e2de99ec5718c00;
    assign coff[6860] = 64'h71d21662c5718c00;
    assign coff[6861] = 64'h2713e35f861c68e4;
    assign coff[6862] = 64'hc5718c008e2de99e;
    assign coff[6863] = 64'h861c68e4d8ec1ca1;
    assign coff[6864] = 64'h6fec5c3bc1e4d0b6;
    assign coff[6865] = 64'h2339db5e84f14ce8;
    assign coff[6866] = 64'hc1e4d0b69013a3c5;
    assign coff[6867] = 64'h84f14ce8dcc624a2;
    assign coff[6868] = 64'h7b0eb318dcc624a2;
    assign coff[6869] = 64'h3e1b2f4a9013a3c5;
    assign coff[6870] = 64'hdcc624a284f14ce8;
    assign coff[6871] = 64'h9013a3c5c1e4d0b6;
    assign coff[6872] = 64'h7f2baf0df173da2b;
    assign coff[6873] = 64'h4fa2f9819bca48fa;
    assign coff[6874] = 64'hf173da2b80d450f3;
    assign coff[6875] = 64'h9bca48fab05d067f;
    assign coff[6876] = 64'h6435b706b05d067f;
    assign coff[6877] = 64'h0e8c25d580d450f3;
    assign coff[6878] = 64'hb05d067f9bca48fa;
    assign coff[6879] = 64'h80d450f3f173da2b;
    assign coff[6880] = 64'h694bffabb738f3a7;
    assign coff[6881] = 64'h16fea10282151709;
    assign coff[6882] = 64'hb738f3a796b40055;
    assign coff[6883] = 64'h82151709e9015efe;
    assign coff[6884] = 64'h7deae8f7e9015efe;
    assign coff[6885] = 64'h48c70c5996b40055;
    assign coff[6886] = 64'he9015efe82151709;
    assign coff[6887] = 64'h96b40055b738f3a7;
    assign coff[6888] = 64'h7d21e393e50ec51d;
    assign coff[6889] = 64'h456e4d4f94778ab1;
    assign coff[6890] = 64'he50ec51d82de1c6d;
    assign coff[6891] = 64'h94778ab1ba91b2b1;
    assign coff[6892] = 64'h6b88754fba91b2b1;
    assign coff[6893] = 64'h1af13ae382de1c6d;
    assign coff[6894] = 64'hba91b2b194778ab1;
    assign coff[6895] = 64'h82de1c6de50ec51d;
    assign coff[6896] = 64'h7578c8b0cd29cbee;
    assign coff[6897] = 64'h2f1e3ced88fce62a;
    assign coff[6898] = 64'hcd29cbee8a873750;
    assign coff[6899] = 64'h88fce62ad0e1c313;
    assign coff[6900] = 64'h770319d6d0e1c313;
    assign coff[6901] = 64'h32d634128a873750;
    assign coff[6902] = 64'hd0e1c31388fce62a;
    assign coff[6903] = 64'h8a873750cd29cbee;
    assign coff[6904] = 64'h7ffbf319fdfccccf;
    assign coff[6905] = 64'h59134f3ea4141672;
    assign coff[6906] = 64'hfdfccccf80040ce7;
    assign coff[6907] = 64'ha4141672a6ecb0c2;
    assign coff[6908] = 64'h5bebe98ea6ecb0c2;
    assign coff[6909] = 64'h0203333180040ce7;
    assign coff[6910] = 64'ha6ecb0c2a4141672;
    assign coff[6911] = 64'h80040ce7fdfccccf;
    assign coff[6912] = 64'h5c660084a76b5c19;
    assign coff[6913] = 64'h02b31961800749e7;
    assign coff[6914] = 64'ha76b5c19a399ff7c;
    assign coff[6915] = 64'h800749e7fd4ce69f;
    assign coff[6916] = 64'h7ff8b619fd4ce69f;
    assign coff[6917] = 64'h5894a3e7a399ff7c;
    assign coff[6918] = 64'hfd4ce69f800749e7;
    assign coff[6919] = 64'ha399ff7ca76b5c19;
    assign coff[6920] = 64'h77436c40d18582ca;
    assign coff[6921] = 64'h3377794b8acd8583;
    assign coff[6922] = 64'hd18582ca88bc93c0;
    assign coff[6923] = 64'h8acd8583cc8886b5;
    assign coff[6924] = 64'h75327a7dcc8886b5;
    assign coff[6925] = 64'h2e7a7d3688bc93c0;
    assign coff[6926] = 64'hcc8886b58acd8583;
    assign coff[6927] = 64'h88bc93c0d18582ca;
    assign coff[6928] = 64'h6be77d74bb25c07d;
    assign coff[6929] = 64'h1b9d1e1a83039a73;
    assign coff[6930] = 64'hbb25c07d9418828c;
    assign coff[6931] = 64'h83039a73e462e1e6;
    assign coff[6932] = 64'h7cfc658de462e1e6;
    assign coff[6933] = 64'h44da3f839418828c;
    assign coff[6934] = 64'he462e1e683039a73;
    assign coff[6935] = 64'h9418828cbb25c07d;
    assign coff[6936] = 64'h7e0a0cd9e9ae85ab;
    assign coff[6937] = 64'h4957810397186b0d;
    assign coff[6938] = 64'he9ae85ab81f5f327;
    assign coff[6939] = 64'h97186b0db6a87efd;
    assign coff[6940] = 64'h68e794f3b6a87efd;
    assign coff[6941] = 64'h16517a5581f5f327;
    assign coff[6942] = 64'hb6a87efd97186b0d;
    assign coff[6943] = 64'h81f5f327e9ae85ab;
    assign coff[6944] = 64'h64a2cd0cb0e70d37;
    assign coff[6945] = 64'h0f3ae1ee80e8c7b0;
    assign coff[6946] = 64'hb0e70d379b5d32f4;
    assign coff[6947] = 64'h80e8c7b0f0c51e12;
    assign coff[6948] = 64'h7f173850f0c51e12;
    assign coff[6949] = 64'h4f18f2c99b5d32f4;
    assign coff[6950] = 64'hf0c51e1280e8c7b0;
    assign coff[6951] = 64'h9b5d32f4b0e70d37;
    assign coff[6952] = 64'h7b3ea95ddd6f687b;
    assign coff[6953] = 64'h3eb4c995906969f8;
    assign coff[6954] = 64'hdd6f687b84c156a3;
    assign coff[6955] = 64'h906969f8c14b366b;
    assign coff[6956] = 64'h6f969608c14b366b;
    assign coff[6957] = 64'h2290978584c156a3;
    assign coff[6958] = 64'hc14b366b906969f8;
    assign coff[6959] = 64'h84c156a3dd6f687b;
    assign coff[6960] = 64'h7222265bc60e33df;
    assign coff[6961] = 64'h27bb45ed865291c4;
    assign coff[6962] = 64'hc60e33df8dddd9a5;
    assign coff[6963] = 64'h865291c4d844ba13;
    assign coff[6964] = 64'h79ad6e3cd844ba13;
    assign coff[6965] = 64'h39f1cc218dddd9a5;
    assign coff[6966] = 64'hd844ba13865291c4;
    assign coff[6967] = 64'h8dddd9a5c60e33df;
    assign coff[6968] = 64'h7f9eb2f8f624a8fa;
    assign coff[6969] = 64'h534566f09eca0e6d;
    assign coff[6970] = 64'hf624a8fa80614d08;
    assign coff[6971] = 64'h9eca0e6dacba9910;
    assign coff[6972] = 64'h6135f193acba9910;
    assign coff[6973] = 64'h09db570680614d08;
    assign coff[6974] = 64'hacba99109eca0e6d;
    assign coff[6975] = 64'h80614d08f624a8fa;
    assign coff[6976] = 64'h60a23322ac0f5256;
    assign coff[6977] = 64'h08f9c2338050a939;
    assign coff[6978] = 64'hac0f52569f5dccde;
    assign coff[6979] = 64'h8050a939f7063dcd;
    assign coff[6980] = 64'h7faf56c7f7063dcd;
    assign coff[6981] = 64'h53f0adaa9f5dccde;
    assign coff[6982] = 64'hf7063dcd8050a939;
    assign coff[6983] = 64'h9f5dccdeac0f5256;
    assign coff[6984] = 64'h79667a44d76df2f6;
    assign coff[6985] = 64'h3927c1558d782694;
    assign coff[6986] = 64'hd76df2f6869985bc;
    assign coff[6987] = 64'h8d782694c6d83eab;
    assign coff[6988] = 64'h7287d96cc6d83eab;
    assign coff[6989] = 64'h28920d0a869985bc;
    assign coff[6990] = 64'hc6d83eab8d782694;
    assign coff[6991] = 64'h869985bcd76df2f6;
    assign coff[6992] = 64'h6f271868c0866767;
    assign coff[6993] = 64'h21b6975f84850271;
    assign coff[6994] = 64'hc086676790d8e798;
    assign coff[6995] = 64'h84850271de4968a1;
    assign coff[6996] = 64'h7b7afd8fde4968a1;
    assign coff[6997] = 64'h3f79989990d8e798;
    assign coff[6998] = 64'hde4968a184850271;
    assign coff[6999] = 64'h90d8e798c0866767;
    assign coff[7000] = 64'h7efb8809efe49fd3;
    assign coff[7001] = 64'h4e66a1059ad20987;
    assign coff[7002] = 64'hefe49fd3810477f7;
    assign coff[7003] = 64'h9ad20987b1995efb;
    assign coff[7004] = 64'h652df679b1995efb;
    assign coff[7005] = 64'h101b602d810477f7;
    assign coff[7006] = 64'hb1995efb9ad20987;
    assign coff[7007] = 64'h810477f7efe49fd3;
    assign coff[7008] = 64'h6865565cb5ef9026;
    assign coff[7009] = 64'h15729d1f81cf477b;
    assign coff[7010] = 64'hb5ef9026979aa9a4;
    assign coff[7011] = 64'h81cf477bea8d62e1;
    assign coff[7012] = 64'h7e30b885ea8d62e1;
    assign coff[7013] = 64'h4a106fda979aa9a4;
    assign coff[7014] = 64'hea8d62e181cf477b;
    assign coff[7015] = 64'h979aa9a4b5ef9026;
    assign coff[7016] = 64'h7ccad656e3862f2a;
    assign coff[7017] = 64'h441b25a8939f7f20;
    assign coff[7018] = 64'he3862f2a833529aa;
    assign coff[7019] = 64'h939f7f20bbe4da58;
    assign coff[7020] = 64'h6c6080e0bbe4da58;
    assign coff[7021] = 64'h1c79d0d6833529aa;
    assign coff[7022] = 64'hbbe4da58939f7f20;
    assign coff[7023] = 64'h833529aae3862f2a;
    assign coff[7024] = 64'h74d6d0b2cbb9bcbb;
    assign coff[7025] = 64'h2da77397886b2bc5;
    assign coff[7026] = 64'hcbb9bcbb8b292f4e;
    assign coff[7027] = 64'h886b2bc5d2588c69;
    assign coff[7028] = 64'h7794d43bd2588c69;
    assign coff[7029] = 64'h344643458b292f4e;
    assign coff[7030] = 64'hd2588c69886b2bc5;
    assign coff[7031] = 64'h8b292f4ecbb9bcbb;
    assign coff[7032] = 64'h7ff32905fc6ac657;
    assign coff[7033] = 64'h57f0d1daa2fe0724;
    assign coff[7034] = 64'hfc6ac657800cd6fb;
    assign coff[7035] = 64'ha2fe0724a80f2e26;
    assign coff[7036] = 64'h5d01f8dca80f2e26;
    assign coff[7037] = 64'h039539a9800cd6fb;
    assign coff[7038] = 64'ha80f2e26a2fe0724;
    assign coff[7039] = 64'h800cd6fbfc6ac657;
    assign coff[7040] = 64'h5e8b63f7a9b6b014;
    assign coff[7041] = 64'h05d6e10c80221db3;
    assign coff[7042] = 64'ha9b6b014a1749c09;
    assign coff[7043] = 64'h80221db3fa291ef4;
    assign coff[7044] = 64'h7fdde24dfa291ef4;
    assign coff[7045] = 64'h56494feca1749c09;
    assign coff[7046] = 64'hfa291ef480221db3;
    assign coff[7047] = 64'ha1749c09a9b6b014;
    assign coff[7048] = 64'h785e3b1cd4765f85;
    assign coff[7049] = 64'h3653cda38c19e669;
    assign coff[7050] = 64'hd4765f8587a1c4e4;
    assign coff[7051] = 64'h8c19e669c9ac325d;
    assign coff[7052] = 64'h73e61997c9ac325d;
    assign coff[7053] = 64'h2b89a07b87a1c4e4;
    assign coff[7054] = 64'hc9ac325d8c19e669;
    assign coff[7055] = 64'h87a1c4e4d4765f85;
    assign coff[7056] = 64'h6d8fbd7abdd0f999;
    assign coff[7057] = 64'h1eac382983bab991;
    assign coff[7058] = 64'hbdd0f99992704286;
    assign coff[7059] = 64'h83bab991e153c7d7;
    assign coff[7060] = 64'h7c45466fe153c7d7;
    assign coff[7061] = 64'h422f066792704286;
    assign coff[7062] = 64'he153c7d783bab991;
    assign coff[7063] = 64'h92704286bdd0f999;
    assign coff[7064] = 64'h7e8c8c4becc81769;
    assign coff[7065] = 64'h4be4eb0898ed47cf;
    assign coff[7066] = 64'hecc81769817373b5;
    assign coff[7067] = 64'h98ed47cfb41b14f8;
    assign coff[7068] = 64'h6712b831b41b14f8;
    assign coff[7069] = 64'h1337e897817373b5;
    assign coff[7070] = 64'hb41b14f898ed47cf;
    assign coff[7071] = 64'h817373b5ecc81769;
    assign coff[7072] = 64'h668bf9cbb36566a8;
    assign coff[7073] = 64'h1258299c8152432c;
    assign coff[7074] = 64'hb36566a899740635;
    assign coff[7075] = 64'h8152432ceda7d664;
    assign coff[7076] = 64'h7eadbcd4eda7d664;
    assign coff[7077] = 64'h4c9a995899740635;
    assign coff[7078] = 64'heda7d6648152432c;
    assign coff[7079] = 64'h99740635b36566a8;
    assign coff[7080] = 64'h7c0e507ee0785d7b;
    assign coff[7081] = 64'h416d030291fbf908;
    assign coff[7082] = 64'he0785d7b83f1af82;
    assign coff[7083] = 64'h91fbf908be92fcfe;
    assign coff[7084] = 64'h6e0406f8be92fcfe;
    assign coff[7085] = 64'h1f87a28583f1af82;
    assign coff[7086] = 64'hbe92fcfe91fbf908;
    assign coff[7087] = 64'h83f1af82e0785d7b;
    assign coff[7088] = 64'h738563b5c8dfb836;
    assign coff[7089] = 64'h2ab4a7b18755910b;
    assign coff[7090] = 64'hc8dfb8368c7a9c4b;
    assign coff[7091] = 64'h8755910bd54b584f;
    assign coff[7092] = 64'h78aa6ef5d54b584f;
    assign coff[7093] = 64'h372047ca8c7a9c4b;
    assign coff[7094] = 64'hd54b584f8755910b;
    assign coff[7095] = 64'h8c7a9c4bc8dfb836;
    assign coff[7096] = 64'h7fd2c900f94732fb;
    assign coff[7097] = 64'h55a1b69da0dcb4ee;
    assign coff[7098] = 64'hf94732fb802d3700;
    assign coff[7099] = 64'ha0dcb4eeaa5e4963;
    assign coff[7100] = 64'h5f234b12aa5e4963;
    assign coff[7101] = 64'h06b8cd05802d3700;
    assign coff[7102] = 64'haa5e4963a0dcb4ee;
    assign coff[7103] = 64'h802d3700f94732fb;
    assign coff[7104] = 64'h62aa1b8dae74e641;
    assign coff[7105] = 64'h0c1b41078092e54a;
    assign coff[7106] = 64'hae74e6419d55e473;
    assign coff[7107] = 64'h8092e54af3e4bef9;
    assign coff[7108] = 64'h7f6d1ab6f3e4bef9;
    assign coff[7109] = 64'h518b19bf9d55e473;
    assign coff[7110] = 64'hf3e4bef98092e54a;
    assign coff[7111] = 64'h9d55e473ae74e641;
    assign coff[7112] = 64'h7a5c00f9da6bc7fa;
    assign coff[7113] = 64'h3bf2e4be8ee81002;
    assign coff[7114] = 64'hda6bc7fa85a3ff07;
    assign coff[7115] = 64'h8ee81002c40d1b42;
    assign coff[7116] = 64'h7117effec40d1b42;
    assign coff[7117] = 64'h2594380685a3ff07;
    assign coff[7118] = 64'hc40d1b428ee81002;
    assign coff[7119] = 64'h85a3ff07da6bc7fa;
    assign coff[7120] = 64'h70ad4f6dc3459ef9;
    assign coff[7121] = 64'h24bbc3b4856255e3;
    assign coff[7122] = 64'hc3459ef98f52b093;
    assign coff[7123] = 64'h856255e3db443c4c;
    assign coff[7124] = 64'h7a9daa1ddb443c4c;
    assign coff[7125] = 64'h3cba61078f52b093;
    assign coff[7126] = 64'hdb443c4c856255e3;
    assign coff[7127] = 64'h8f52b093c3459ef9;
    assign coff[7128] = 64'h7f56eef5f303a416;
    assign coff[7129] = 64'h50dc40059cc66573;
    assign coff[7130] = 64'hf303a41680a9110b;
    assign coff[7131] = 64'h9cc66573af23bffb;
    assign coff[7132] = 64'h63399a8daf23bffb;
    assign coff[7133] = 64'h0cfc5bea80a9110b;
    assign coff[7134] = 64'haf23bffb9cc66573;
    assign coff[7135] = 64'h80a9110bf303a416;
    assign coff[7136] = 64'h6a2e99c0b885256f;
    assign coff[7137] = 64'h1889c1f3825fc155;
    assign coff[7138] = 64'hb885256f95d16640;
    assign coff[7139] = 64'h825fc155e7763e0d;
    assign coff[7140] = 64'h7da03eabe7763e0d;
    assign coff[7141] = 64'h477ada9195d16640;
    assign coff[7142] = 64'he7763e0d825fc155;
    assign coff[7143] = 64'h95d16640b885256f;
    assign coff[7144] = 64'h7d741dd2e69864f9;
    assign coff[7145] = 64'h46bec7b89553bb8e;
    assign coff[7146] = 64'he69864f9828be22e;
    assign coff[7147] = 64'h9553bb8eb9413848;
    assign coff[7148] = 64'h6aac4472b9413848;
    assign coff[7149] = 64'h19679b07828be22e;
    assign coff[7150] = 64'hb94138489553bb8e;
    assign coff[7151] = 64'h828be22ee69864f9;
    assign coff[7152] = 64'h7616394cce9bd0dd;
    assign coff[7153] = 64'h3093353a89933725;
    assign coff[7154] = 64'hce9bd0dd89e9c6b4;
    assign coff[7155] = 64'h89933725cf6ccac6;
    assign coff[7156] = 64'h766cc8dbcf6ccac6;
    assign coff[7157] = 64'h31642f2389e9c6b4;
    assign coff[7158] = 64'hcf6ccac689933725;
    assign coff[7159] = 64'h89e9c6b4ce9bd0dd;
    assign coff[7160] = 64'h7fffce09ff8ee724;
    assign coff[7161] = 64'h5a325d82a52db0f7;
    assign coff[7162] = 64'hff8ee724800031f7;
    assign coff[7163] = 64'ha52db0f7a5cda27e;
    assign coff[7164] = 64'h5ad24f09a5cda27e;
    assign coff[7165] = 64'h007118dc800031f7;
    assign coff[7166] = 64'ha5cda27ea52db0f7;
    assign coff[7167] = 64'h800031f7ff8ee724;
    assign coff[7168] = 64'h5b07609da60331b1;
    assign coff[7169] = 64'h00bc7e9980008aca;
    assign coff[7170] = 64'ha60331b1a4f89f63;
    assign coff[7171] = 64'h80008acaff438167;
    assign coff[7172] = 64'h7fff7536ff438167;
    assign coff[7173] = 64'h59fcce4fa4f89f63;
    assign coff[7174] = 64'hff43816780008aca;
    assign coff[7175] = 64'ha4f89f63a60331b1;
    assign coff[7176] = 64'h7689513fcfb2953f;
    assign coff[7177] = 64'h31a9b5a08a06f339;
    assign coff[7178] = 64'hcfb2953f8976aec1;
    assign coff[7179] = 64'h8a06f339ce564a60;
    assign coff[7180] = 64'h75f90cc7ce564a60;
    assign coff[7181] = 64'h304d6ac18976aec1;
    assign coff[7182] = 64'hce564a608a06f339;
    assign coff[7183] = 64'h8976aec1cfb2953f;
    assign coff[7184] = 64'h6ad5de0fb9801a70;
    assign coff[7185] = 64'h19b17c8f829aeee1;
    assign coff[7186] = 64'hb9801a70952a21f1;
    assign coff[7187] = 64'h829aeee1e64e8371;
    assign coff[7188] = 64'h7d65111fe64e8371;
    assign coff[7189] = 64'h467fe590952a21f1;
    assign coff[7190] = 64'he64e8371829aeee1;
    assign coff[7191] = 64'h952a21f1b9801a70;
    assign coff[7192] = 64'h7dae9d21e7c0423d;
    assign coff[7193] = 64'h47b95a0695fb9394;
    assign coff[7194] = 64'he7c0423d825162df;
    assign coff[7195] = 64'h95fb9394b846a5fa;
    assign coff[7196] = 64'h6a046c6cb846a5fa;
    assign coff[7197] = 64'h183fbdc3825162df;
    assign coff[7198] = 64'hb846a5fa95fb9394;
    assign coff[7199] = 64'h825162dfe7c0423d;
    assign coff[7200] = 64'h63692ac7af5e40c7;
    assign coff[7201] = 64'h0d475c0080b0cd57;
    assign coff[7202] = 64'haf5e40c79c96d539;
    assign coff[7203] = 64'h80b0cd57f2b8a400;
    assign coff[7204] = 64'h7f4f32a9f2b8a400;
    assign coff[7205] = 64'h50a1bf399c96d539;
    assign coff[7206] = 64'hf2b8a40080b0cd57;
    assign coff[7207] = 64'h9c96d539af5e40c7;
    assign coff[7208] = 64'h7ab3381ddb8c7cb1;
    assign coff[7209] = 64'h3cfcb5c48f7689b0;
    assign coff[7210] = 64'hdb8c7cb1854cc7e3;
    assign coff[7211] = 64'h8f7689b0c3034a3c;
    assign coff[7212] = 64'h70897650c3034a3c;
    assign coff[7213] = 64'h2473834f854cc7e3;
    assign coff[7214] = 64'hc3034a3c8f7689b0;
    assign coff[7215] = 64'h854cc7e3db8c7cb1;
    assign coff[7216] = 64'h713b2c6ec44fc3be;
    assign coff[7217] = 64'h25dc44d985ba3707;
    assign coff[7218] = 64'hc44fc3be8ec4d392;
    assign coff[7219] = 64'h85ba3707da23bb27;
    assign coff[7220] = 64'h7a45c8f9da23bb27;
    assign coff[7221] = 64'h3bb03c428ec4d392;
    assign coff[7222] = 64'hda23bb2785ba3707;
    assign coff[7223] = 64'h8ec4d392c44fc3be;
    assign coff[7224] = 64'h7f742637f42fd079;
    assign coff[7225] = 64'h51c529d79d85fe02;
    assign coff[7226] = 64'hf42fd079808bd9c9;
    assign coff[7227] = 64'h9d85fe02ae3ad629;
    assign coff[7228] = 64'h627a01feae3ad629;
    assign coff[7229] = 64'h0bd02f87808bd9c9;
    assign coff[7230] = 64'hae3ad6299d85fe02;
    assign coff[7231] = 64'h808bd9c9f42fd079;
    assign coff[7232] = 64'h5f55ab82aa9662af;
    assign coff[7233] = 64'h07041726803142cf;
    assign coff[7234] = 64'haa9662afa0aa547e;
    assign coff[7235] = 64'h803142cff8fbe8da;
    assign coff[7236] = 64'h7fcebd31f8fbe8da;
    assign coff[7237] = 64'h55699d51a0aa547e;
    assign coff[7238] = 64'hf8fbe8da803142cf;
    assign coff[7239] = 64'ha0aa547eaa9662af;
    assign coff[7240] = 64'h78c381e2d59273ab;
    assign coff[7241] = 64'h37644a608c9b2926;
    assign coff[7242] = 64'hd59273ab873c7e1e;
    assign coff[7243] = 64'h8c9b2926c89bb5a0;
    assign coff[7244] = 64'h7364d6dac89bb5a0;
    assign coff[7245] = 64'h2a6d8c55873c7e1e;
    assign coff[7246] = 64'hc89bb5a08c9b2926;
    assign coff[7247] = 64'h873c7e1ed59273ab;
    assign coff[7248] = 64'h6e2a7ddbbed3d64f;
    assign coff[7249] = 64'h1fd0b03a8404579d;
    assign coff[7250] = 64'hbed3d64f91d58225;
    assign coff[7251] = 64'h8404579de02f4fc6;
    assign coff[7252] = 64'h7bfba863e02f4fc6;
    assign coff[7253] = 64'h412c29b191d58225;
    assign coff[7254] = 64'he02f4fc68404579d;
    assign coff[7255] = 64'h91d58225bed3d64f;
    assign coff[7256] = 64'h7eb8751eedf2783f;
    assign coff[7257] = 64'h4cd6f3bb99a13795;
    assign coff[7258] = 64'hedf2783f81478ae2;
    assign coff[7259] = 64'h99a13795b3290c45;
    assign coff[7260] = 64'h665ec86bb3290c45;
    assign coff[7261] = 64'h120d87c181478ae2;
    assign coff[7262] = 64'hb3290c4599a13795;
    assign coff[7263] = 64'h81478ae2edf2783f;
    assign coff[7264] = 64'h673f5ae0b457d92f;
    assign coff[7265] = 64'h13827062817edbb9;
    assign coff[7266] = 64'hb457d92f98c0a520;
    assign coff[7267] = 64'h817edbb9ec7d8f9e;
    assign coff[7268] = 64'h7e812447ec7d8f9e;
    assign coff[7269] = 64'h4ba826d198c0a520;
    assign coff[7270] = 64'hec7d8f9e817edbb9;
    assign coff[7271] = 64'h98c0a520b457d92f;
    assign coff[7272] = 64'h7c574236e19d00b6;
    assign coff[7273] = 64'h426f8463929751c9;
    assign coff[7274] = 64'he19d00b683a8bdca;
    assign coff[7275] = 64'h929751c9bd907b9d;
    assign coff[7276] = 64'h6d68ae37bd907b9d;
    assign coff[7277] = 64'h1e62ff4a83a8bdca;
    assign coff[7278] = 64'hbd907b9d929751c9;
    assign coff[7279] = 64'h83a8bdcae19d00b6;
    assign coff[7280] = 64'h740605d9c9f080e7;
    assign coff[7281] = 64'h2bd07ffe87bb7f16;
    assign coff[7282] = 64'hc9f080e78bf9fa27;
    assign coff[7283] = 64'h87bb7f16d42f8002;
    assign coff[7284] = 64'h784480ead42f8002;
    assign coff[7285] = 64'h360f7f198bf9fa27;
    assign coff[7286] = 64'hd42f800287bb7f16;
    assign coff[7287] = 64'h8bf9fa27c9f080e7;
    assign coff[7288] = 64'h7fe13cacfa7471cc;
    assign coff[7289] = 64'h5680f1eaa1a7801b;
    assign coff[7290] = 64'hfa7471cc801ec354;
    assign coff[7291] = 64'ha1a7801ba97f0e16;
    assign coff[7292] = 64'h5e587fe5a97f0e16;
    assign coff[7293] = 64'h058b8e34801ec354;
    assign coff[7294] = 64'ha97f0e16a1a7801b;
    assign coff[7295] = 64'h801ec354fa7471cc;
    assign coff[7296] = 64'h5d35b5dba84606a0;
    assign coff[7297] = 64'h03e09767800f0978;
    assign coff[7298] = 64'ha84606a0a2ca4a25;
    assign coff[7299] = 64'h800f0978fc1f6899;
    assign coff[7300] = 64'h7ff0f688fc1f6899;
    assign coff[7301] = 64'h57b9f960a2ca4a25;
    assign coff[7302] = 64'hfc1f6899800f0978;
    assign coff[7303] = 64'ha2ca4a25a84606a0;
    assign coff[7304] = 64'h77afa3f5d29f04c2;
    assign coff[7305] = 64'h348b0d1c8b480e5f;
    assign coff[7306] = 64'hd29f04c288505c0b;
    assign coff[7307] = 64'h8b480e5fcb74f2e4;
    assign coff[7308] = 64'h74b7f1a1cb74f2e4;
    assign coff[7309] = 64'h2d60fb3e88505c0b;
    assign coff[7310] = 64'hcb74f2e48b480e5f;
    assign coff[7311] = 64'h88505c0bd29f04c2;
    assign coff[7312] = 64'h6c888c36bc24bd02;
    assign coff[7313] = 64'h1cc34e1f8346055e;
    assign coff[7314] = 64'hbc24bd02937773ca;
    assign coff[7315] = 64'h8346055ee33cb1e1;
    assign coff[7316] = 64'h7cb9faa2e33cb1e1;
    assign coff[7317] = 64'h43db42fe937773ca;
    assign coff[7318] = 64'he33cb1e18346055e;
    assign coff[7319] = 64'h937773cabc24bd02;
    assign coff[7320] = 64'h7e3d44ddead7bba3;
    assign coff[7321] = 64'h4a4de18297c65c5c;
    assign coff[7322] = 64'head7bba381c2bb23;
    assign coff[7323] = 64'h97c65c5cb5b21e7e;
    assign coff[7324] = 64'h6839a3a4b5b21e7e;
    assign coff[7325] = 64'h1528445d81c2bb23;
    assign coff[7326] = 64'hb5b21e7e97c65c5c;
    assign coff[7327] = 64'h81c2bb23ead7bba3;
    assign coff[7328] = 64'h655c137db1d50616;
    assign coff[7329] = 64'h106629e1810e0adc;
    assign coff[7330] = 64'hb1d506169aa3ec83;
    assign coff[7331] = 64'h810e0adcef99d61f;
    assign coff[7332] = 64'h7ef1f524ef99d61f;
    assign coff[7333] = 64'h4e2af9ea9aa3ec83;
    assign coff[7334] = 64'hef99d61f810e0adc;
    assign coff[7335] = 64'h9aa3ec83b1d50616;
    assign coff[7336] = 64'h7b8ec3f8de922adf;
    assign coff[7337] = 64'h3fbb070290fe5eab;
    assign coff[7338] = 64'hde922adf84713c08;
    assign coff[7339] = 64'h90fe5eabc044f8fe;
    assign coff[7340] = 64'h6f01a155c044f8fe;
    assign coff[7341] = 64'h216dd52184713c08;
    assign coff[7342] = 64'hc044f8fe90fe5eab;
    assign coff[7343] = 64'h84713c08de922adf;
    assign coff[7344] = 64'h72a9705cc71bbf62;
    assign coff[7345] = 64'h28d988b886b180ae;
    assign coff[7346] = 64'hc71bbf628d568fa4;
    assign coff[7347] = 64'h86b180aed7267748;
    assign coff[7348] = 64'h794e7f52d7267748;
    assign coff[7349] = 64'h38e4409e8d568fa4;
    assign coff[7350] = 64'hd726774886b180ae;
    assign coff[7351] = 64'h8d568fa4c71bbf62;
    assign coff[7352] = 64'h7fb48a1ef75175c6;
    assign coff[7353] = 64'h54298b179f8f4f80;
    assign coff[7354] = 64'hf75175c6804b75e2;
    assign coff[7355] = 64'h9f8f4f80abd674e9;
    assign coff[7356] = 64'h6070b080abd674e9;
    assign coff[7357] = 64'h08ae8a3a804b75e2;
    assign coff[7358] = 64'habd674e99f8f4f80;
    assign coff[7359] = 64'h804b75e2f75175c6;
    assign coff[7360] = 64'h6166edb0acf3ea87;
    assign coff[7361] = 64'h0a2681ed8067318a;
    assign coff[7362] = 64'hacf3ea879e991250;
    assign coff[7363] = 64'h8067318af5d97e13;
    assign coff[7364] = 64'h7f98ce76f5d97e13;
    assign coff[7365] = 64'h530c15799e991250;
    assign coff[7366] = 64'hf5d97e138067318a;
    assign coff[7367] = 64'h9e991250acf3ea87;
    assign coff[7368] = 64'h79c4c07ed88c6d7b;
    assign coff[7369] = 64'h3a34fcf98e000f44;
    assign coff[7370] = 64'hd88c6d7b863b3f82;
    assign coff[7371] = 64'h8e000f44c5cb0307;
    assign coff[7372] = 64'h71fff0bcc5cb0307;
    assign coff[7373] = 64'h27739285863b3f82;
    assign coff[7374] = 64'hc5cb03078e000f44;
    assign coff[7375] = 64'h863b3f82d88c6d7b;
    assign coff[7376] = 64'h6fbb728ac18cfc63;
    assign coff[7377] = 64'h22d92a6184d5c844;
    assign coff[7378] = 64'hc18cfc6390448d76;
    assign coff[7379] = 64'h84d5c844dd26d59f;
    assign coff[7380] = 64'h7b2a37bcdd26d59f;
    assign coff[7381] = 64'h3e73039d90448d76;
    assign coff[7382] = 64'hdd26d59f84d5c844;
    assign coff[7383] = 64'h90448d76c18cfc63;
    assign coff[7384] = 64'h7f201ae5f10ffd85;
    assign coff[7385] = 64'h4f542c989b8bdc05;
    assign coff[7386] = 64'hf10ffd8580dfe51b;
    assign coff[7387] = 64'h9b8bdc05b0abd368;
    assign coff[7388] = 64'h647423fbb0abd368;
    assign coff[7389] = 64'h0ef0027b80dfe51b;
    assign coff[7390] = 64'hb0abd3689b8bdc05;
    assign coff[7391] = 64'h80dfe51bf10ffd85;
    assign coff[7392] = 64'h6912b66cb6e656f1;
    assign coff[7393] = 64'h169bb4b782032e88;
    assign coff[7394] = 64'hb6e656f196ed4994;
    assign coff[7395] = 64'h82032e88e9644b49;
    assign coff[7396] = 64'h7dfcd178e9644b49;
    assign coff[7397] = 64'h4919a90f96ed4994;
    assign coff[7398] = 64'he9644b4982032e88;
    assign coff[7399] = 64'h96ed4994b6e656f1;
    assign coff[7400] = 64'h7d0c93ebe4ac861b;
    assign coff[7401] = 64'h4519c321944123fa;
    assign coff[7402] = 64'he4ac861b82f36c15;
    assign coff[7403] = 64'h944123fabae63cdf;
    assign coff[7404] = 64'h6bbedc06bae63cdf;
    assign coff[7405] = 64'h1b5379e582f36c15;
    assign coff[7406] = 64'hbae63cdf944123fa;
    assign coff[7407] = 64'h82f36c15e4ac861b;
    assign coff[7408] = 64'h7550b725cccd988a;
    assign coff[7409] = 64'h2ec0b5a088d8093a;
    assign coff[7410] = 64'hcccd988a8aaf48db;
    assign coff[7411] = 64'h88d8093ad13f4a60;
    assign coff[7412] = 64'h7727f6c6d13f4a60;
    assign coff[7413] = 64'h333267768aaf48db;
    assign coff[7414] = 64'hd13f4a6088d8093a;
    assign coff[7415] = 64'h8aaf48dbcccd988a;
    assign coff[7416] = 64'h7ffa36fcfd9848b9;
    assign coff[7417] = 64'h58cb01e1a3ce3d25;
    assign coff[7418] = 64'hfd9848b98005c904;
    assign coff[7419] = 64'ha3ce3d25a734fe1f;
    assign coff[7420] = 64'h5c31c2dba734fe1f;
    assign coff[7421] = 64'h0267b7478005c904;
    assign coff[7422] = 64'ha734fe1fa3ce3d25;
    assign coff[7423] = 64'h8005c904fd9848b9;
    assign coff[7424] = 64'h5c2051dba722e5a3;
    assign coff[7425] = 64'h024e966280055296;
    assign coff[7426] = 64'ha722e5a3a3dfae25;
    assign coff[7427] = 64'h80055296fdb1699e;
    assign coff[7428] = 64'h7ffaad6afdb1699e;
    assign coff[7429] = 64'h58dd1a5da3dfae25;
    assign coff[7430] = 64'hfdb1699e80055296;
    assign coff[7431] = 64'ha3dfae25a722e5a3;
    assign coff[7432] = 64'h771ec66ed127e5d7;
    assign coff[7433] = 64'h331b5d918aa53daf;
    assign coff[7434] = 64'hd127e5d788e13992;
    assign coff[7435] = 64'h8aa53dafcce4a26f;
    assign coff[7436] = 64'h755ac251cce4a26f;
    assign coff[7437] = 64'h2ed81a2988e13992;
    assign coff[7438] = 64'hcce4a26f8aa53daf;
    assign coff[7439] = 64'h88e13992d127e5d7;
    assign coff[7440] = 64'h6bb14892bad11652;
    assign coff[7441] = 64'h1b3aebb682ee10ef;
    assign coff[7442] = 64'hbad11652944eb76e;
    assign coff[7443] = 64'h82ee10efe4c5144a;
    assign coff[7444] = 64'h7d11ef11e4c5144a;
    assign coff[7445] = 64'h452ee9ae944eb76e;
    assign coff[7446] = 64'he4c5144a82ee10ef;
    assign coff[7447] = 64'h944eb76ebad11652;
    assign coff[7448] = 64'h7df85ea0e94b8ee5;
    assign coff[7449] = 64'h4905061a96def12f;
    assign coff[7450] = 64'he94b8ee58207a160;
    assign coff[7451] = 64'h96def12fb6faf9e6;
    assign coff[7452] = 64'h69210ed1b6faf9e6;
    assign coff[7453] = 64'h16b4711b8207a160;
    assign coff[7454] = 64'hb6faf9e696def12f;
    assign coff[7455] = 64'h8207a160e94b8ee5;
    assign coff[7456] = 64'h64648e8cb0981b96;
    assign coff[7457] = 64'h0ed70c2c80dcf8b7;
    assign coff[7458] = 64'hb0981b969b9b7174;
    assign coff[7459] = 64'h80dcf8b7f128f3d4;
    assign coff[7460] = 64'h7f230749f128f3d4;
    assign coff[7461] = 64'h4f67e46a9b9b7174;
    assign coff[7462] = 64'hf128f3d480dcf8b7;
    assign coff[7463] = 64'h9b9b7174b0981b96;
    assign coff[7464] = 64'h7b235db2dd0ea759;
    assign coff[7465] = 64'h3e5d122290384c93;
    assign coff[7466] = 64'hdd0ea75984dca24e;
    assign coff[7467] = 64'h90384c93c1a2edde;
    assign coff[7468] = 64'h6fc7b36dc1a2edde;
    assign coff[7469] = 64'h22f158a784dca24e;
    assign coff[7470] = 64'hc1a2edde90384c93;
    assign coff[7471] = 64'h84dca24edd0ea759;
    assign coff[7472] = 64'h71f480bcc5b4a1e5;
    assign coff[7473] = 64'h275ba901863382cf;
    assign coff[7474] = 64'hc5b4a1e58e0b7f44;
    assign coff[7475] = 64'h863382cfd8a456ff;
    assign coff[7476] = 64'h79cc7d31d8a456ff;
    assign coff[7477] = 64'h3a4b5e1b8e0b7f44;
    assign coff[7478] = 64'hd8a456ff863382cf;
    assign coff[7479] = 64'h8e0b7f44c5b4a1e5;
    assign coff[7480] = 64'h7f96cdc9f5c0708d;
    assign coff[7481] = 64'h52f8f3e99e88c5c9;
    assign coff[7482] = 64'hf5c0708d80693237;
    assign coff[7483] = 64'h9e88c5c9ad070c17;
    assign coff[7484] = 64'h61773a37ad070c17;
    assign coff[7485] = 64'h0a3f8f7380693237;
    assign coff[7486] = 64'had070c179e88c5c9;
    assign coff[7487] = 64'h80693237f5c0708d;
    assign coff[7488] = 64'h6060282fabc386ec;
    assign coff[7489] = 64'h089576e58049c3f3;
    assign coff[7490] = 64'habc386ec9f9fd7d1;
    assign coff[7491] = 64'h8049c3f3f76a891b;
    assign coff[7492] = 64'h7fb63c0df76a891b;
    assign coff[7493] = 64'h543c79149f9fd7d1;
    assign coff[7494] = 64'hf76a891b8049c3f3;
    assign coff[7495] = 64'h9f9fd7d1abc386ec;
    assign coff[7496] = 64'h794677a6d70ea688;
    assign coff[7497] = 64'h38cdbbfc8d4b662a;
    assign coff[7498] = 64'hd70ea68886b9885a;
    assign coff[7499] = 64'h8d4b662ac7324404;
    assign coff[7500] = 64'h72b499d6c7324404;
    assign coff[7501] = 64'h28f1597886b9885a;
    assign coff[7502] = 64'hc73244048d4b662a;
    assign coff[7503] = 64'h86b9885ad70ea688;
    assign coff[7504] = 64'h6ef51bbec02f2e6f;
    assign coff[7505] = 64'h215591cc846aae16;
    assign coff[7506] = 64'hc02f2e6f910ae442;
    assign coff[7507] = 64'h846aae16deaa6e34;
    assign coff[7508] = 64'h7b9551eadeaa6e34;
    assign coff[7509] = 64'h3fd0d191910ae442;
    assign coff[7510] = 64'hdeaa6e34846aae16;
    assign coff[7511] = 64'h910ae442c02f2e6f;
    assign coff[7512] = 64'h7eeeba62ef80e97a;
    assign coff[7513] = 64'h4e1711849a949552;
    assign coff[7514] = 64'hef80e97a8111459e;
    assign coff[7515] = 64'h9a949552b1e8ee7c;
    assign coff[7516] = 64'h656b6aaeb1e8ee7c;
    assign coff[7517] = 64'h107f16868111459e;
    assign coff[7518] = 64'hb1e8ee7c9a949552;
    assign coff[7519] = 64'h8111459eef80e97a;
    assign coff[7520] = 64'h682b0ab1b59da8ff;
    assign coff[7521] = 64'h150f7a7a81be9617;
    assign coff[7522] = 64'hb59da8ff97d4f54f;
    assign coff[7523] = 64'h81be9617eaf08586;
    assign coff[7524] = 64'h7e4169e9eaf08586;
    assign coff[7525] = 64'h4a62570197d4f54f;
    assign coff[7526] = 64'heaf0858681be9617;
    assign coff[7527] = 64'h97d4f54fb59da8ff;
    assign coff[7528] = 64'h7cb45272e3243500;
    assign coff[7529] = 64'h43c5f234936a230a;
    assign coff[7530] = 64'he3243500834bad8e;
    assign coff[7531] = 64'h936a230abc3a0dcc;
    assign coff[7532] = 64'h6c95dcf6bc3a0dcc;
    assign coff[7533] = 64'h1cdbcb00834bad8e;
    assign coff[7534] = 64'hbc3a0dcc936a230a;
    assign coff[7535] = 64'h834bad8ee3243500;
    assign coff[7536] = 64'h74ad9e46cb5e08fe;
    assign coff[7537] = 64'h2d497a4a8847755d;
    assign coff[7538] = 64'hcb5e08fe8b5261ba;
    assign coff[7539] = 64'h8847755dd2b685b6;
    assign coff[7540] = 64'h77b88aa3d2b685b6;
    assign coff[7541] = 64'h34a1f7028b5261ba;
    assign coff[7542] = 64'hd2b685b68847755d;
    assign coff[7543] = 64'h8b5261bacb5e08fe;
    assign coff[7544] = 64'h7ff0312cfc0649a5;
    assign coff[7545] = 64'h57a7aa73a2b91254;
    assign coff[7546] = 64'hfc0649a5800fced4;
    assign coff[7547] = 64'ha2b91254a858558d;
    assign coff[7548] = 64'h5d46edaca858558d;
    assign coff[7549] = 64'h03f9b65b800fced4;
    assign coff[7550] = 64'ha858558da2b91254;
    assign coff[7551] = 64'h800fced4fc0649a5;
    assign coff[7552] = 64'h5e4781eda96c896c;
    assign coff[7553] = 64'h05727228801daf11;
    assign coff[7554] = 64'ha96c896ca1b87e13;
    assign coff[7555] = 64'h801daf11fa8d8dd8;
    assign coff[7556] = 64'h7fe250effa8d8dd8;
    assign coff[7557] = 64'h56937694a1b87e13;
    assign coff[7558] = 64'hfa8d8dd8801daf11;
    assign coff[7559] = 64'ha1b87e13a96c896c;
    assign coff[7560] = 64'h783be43ed417e38c;
    assign coff[7561] = 64'h35f8b6148bef5f02;
    assign coff[7562] = 64'hd417e38c87c41bc2;
    assign coff[7563] = 64'h8bef5f02ca0749ec;
    assign coff[7564] = 64'h7410a0feca0749ec;
    assign coff[7565] = 64'h2be81c7487c41bc2;
    assign coff[7566] = 64'hca0749ec8bef5f02;
    assign coff[7567] = 64'h87c41bc2d417e38c;
    assign coff[7568] = 64'h6d5ba0b0bd7b0167;
    assign coff[7569] = 64'h1e4a94a783a2c8c9;
    assign coff[7570] = 64'hbd7b016792a45f50;
    assign coff[7571] = 64'h83a2c8c9e1b56b59;
    assign coff[7572] = 64'h7c5d3737e1b56b59;
    assign coff[7573] = 64'h4284fe9992a45f50;
    assign coff[7574] = 64'he1b56b5983a2c8c9;
    assign coff[7575] = 64'h92a45f50bd7b0167;
    assign coff[7576] = 64'h7e7d4d2fec64b930;
    assign coff[7577] = 64'h4b93df9398b1cc30;
    assign coff[7578] = 64'hec64b9308182b2d1;
    assign coff[7579] = 64'h98b1cc30b46c206d;
    assign coff[7580] = 64'h674e33d0b46c206d;
    assign coff[7581] = 64'h139b46d08182b2d1;
    assign coff[7582] = 64'hb46c206d98b1cc30;
    assign coff[7583] = 64'h8182b2d1ec64b930;
    assign coff[7584] = 64'h664fb010b314f410;
    assign coff[7585] = 64'h11f4a5bd814401e4;
    assign coff[7586] = 64'hb314f41099b04ff0;
    assign coff[7587] = 64'h814401e4ee0b5a43;
    assign coff[7588] = 64'h7ebbfe1cee0b5a43;
    assign coff[7589] = 64'h4ceb0bf099b04ff0;
    assign coff[7590] = 64'hee0b5a43814401e4;
    assign coff[7591] = 64'h99b04ff0b314f410;
    assign coff[7592] = 64'h7bf566cbe016f852;
    assign coff[7593] = 64'h411686e491c8b857;
    assign coff[7594] = 64'he016f852840a9935;
    assign coff[7595] = 64'h91c8b857bee9791c;
    assign coff[7596] = 64'h6e3747a9bee9791c;
    assign coff[7597] = 64'h1fe907ae840a9935;
    assign coff[7598] = 64'hbee9791c91c8b857;
    assign coff[7599] = 64'h840a9935e016f852;
    assign coff[7600] = 64'h7359f456c8850e5d;
    assign coff[7601] = 64'h2a55d54587342bc9;
    assign coff[7602] = 64'hc8850e5d8ca60baa;
    assign coff[7603] = 64'h87342bc9d5aa2abb;
    assign coff[7604] = 64'h78cbd437d5aa2abb;
    assign coff[7605] = 64'h377af1a38ca60baa;
    assign coff[7606] = 64'hd5aa2abb87342bc9;
    assign coff[7607] = 64'h8ca60baac8850e5d;
    assign coff[7608] = 64'h7fcd5a11f8e2d0ae;
    assign coff[7609] = 64'h5556e3a1a0999107;
    assign coff[7610] = 64'hf8e2d0ae8032a5ef;
    assign coff[7611] = 64'ha0999107aaa91c5f;
    assign coff[7612] = 64'h5f666ef9aaa91c5f;
    assign coff[7613] = 64'h071d2f528032a5ef;
    assign coff[7614] = 64'haaa91c5fa0999107;
    assign coff[7615] = 64'h8032a5eff8e2d0ae;
    assign coff[7616] = 64'h6269f1e1ae2781c4;
    assign coff[7617] = 64'h0bb728c780898a72;
    assign coff[7618] = 64'hae2781c49d960e1f;
    assign coff[7619] = 64'h80898a72f448d739;
    assign coff[7620] = 64'h7f76758ef448d739;
    assign coff[7621] = 64'h51d87e3c9d960e1f;
    assign coff[7622] = 64'hf448d73980898a72;
    assign coff[7623] = 64'h9d960e1fae2781c4;
    assign coff[7624] = 64'h7a3e578bda0bb9cb;
    assign coff[7625] = 64'h3b99ff7d8eb91d7c;
    assign coff[7626] = 64'hda0bb9cb85c1a875;
    assign coff[7627] = 64'h8eb91d7cc4660083;
    assign coff[7628] = 64'h7146e284c4660083;
    assign coff[7629] = 64'h25f4463585c1a875;
    assign coff[7630] = 64'hc46600838eb91d7c;
    assign coff[7631] = 64'h85c1a875da0bb9cb;
    assign coff[7632] = 64'h707d7a98c2ed32af;
    assign coff[7633] = 64'h245b6b078545a204;
    assign coff[7634] = 64'hc2ed32af8f828568;
    assign coff[7635] = 64'h8545a204dba494f9;
    assign coff[7636] = 64'h7aba5dfcdba494f9;
    assign coff[7637] = 64'h3d12cd518f828568;
    assign coff[7638] = 64'hdba494f98545a204;
    assign coff[7639] = 64'h8f828568c2ed32af;
    assign coff[7640] = 64'h7f4c94bef29fa4fd;
    assign coff[7641] = 64'h508e38bd9c870224;
    assign coff[7642] = 64'hf29fa4fd80b36b42;
    assign coff[7643] = 64'h9c870224af71c743;
    assign coff[7644] = 64'h6378fddcaf71c743;
    assign coff[7645] = 64'h0d605b0380b36b42;
    assign coff[7646] = 64'haf71c7439c870224;
    assign coff[7647] = 64'h80b36b42f29fa4fd;
    assign coff[7648] = 64'h69f65523b831d659;
    assign coff[7649] = 64'h18270fd3824ca268;
    assign coff[7650] = 64'hb831d6599609aadd;
    assign coff[7651] = 64'h824ca268e7d8f02d;
    assign coff[7652] = 64'h7db35d98e7d8f02d;
    assign coff[7653] = 64'h47ce29a79609aadd;
    assign coff[7654] = 64'he7d8f02d824ca268;
    assign coff[7655] = 64'h9609aaddb831d659;
    assign coff[7656] = 64'h7d600338e635e4e9;
    assign coff[7657] = 64'h466aea12951c4c4e;
    assign coff[7658] = 64'he635e4e9829ffcc8;
    assign coff[7659] = 64'h951c4c4eb99515ee;
    assign coff[7660] = 64'h6ae3b3b2b99515ee;
    assign coff[7661] = 64'h19ca1b17829ffcc8;
    assign coff[7662] = 64'hb99515ee951c4c4e;
    assign coff[7663] = 64'h829ffcc8e635e4e9;
    assign coff[7664] = 64'h75ef4a2cce3f215f;
    assign coff[7665] = 64'h30362389896d3518;
    assign coff[7666] = 64'hce3f215f8a10b5d4;
    assign coff[7667] = 64'h896d3518cfc9dc77;
    assign coff[7668] = 64'h7692cae8cfc9dc77;
    assign coff[7669] = 64'h31c0dea18a10b5d4;
    assign coff[7670] = 64'hcfc9dc77896d3518;
    assign coff[7671] = 64'h8a10b5d4ce3f215f;
    assign coff[7672] = 64'h7fff4dbbff2a5f8b;
    assign coff[7673] = 64'h59eaecf8a4e6f5e0;
    assign coff[7674] = 64'hff2a5f8b8000b245;
    assign coff[7675] = 64'ha4e6f5e0a6151308;
    assign coff[7676] = 64'h5b190a20a6151308;
    assign coff[7677] = 64'h00d5a0758000b245;
    assign coff[7678] = 64'ha6151308a4e6f5e0;
    assign coff[7679] = 64'h8000b245ff2a5f8b;
    assign coff[7680] = 64'h5b944a37a6929d57;
    assign coff[7681] = 64'h01858c5e800250c9;
    assign coff[7682] = 64'ha6929d57a46bb5c9;
    assign coff[7683] = 64'h800250c9fe7a73a2;
    assign coff[7684] = 64'h7ffdaf37fe7a73a2;
    assign coff[7685] = 64'h596d62a9a46bb5c9;
    assign coff[7686] = 64'hfe7a73a2800250c9;
    assign coff[7687] = 64'ha46bb5c9a6929d57;
    assign coff[7688] = 64'h76d49e70d06d02da;
    assign coff[7689] = 64'h3262c7c18a55874a;
    assign coff[7690] = 64'hd06d02da892b6190;
    assign coff[7691] = 64'h8a55874acd9d383f;
    assign coff[7692] = 64'h75aa78b6cd9d383f;
    assign coff[7693] = 64'h2f92fd26892b6190;
    assign coff[7694] = 64'hcd9d383f8a55874a;
    assign coff[7695] = 64'h892b6190d06d02da;
    assign coff[7696] = 64'h6b4417a6ba284237;
    assign coff[7697] = 64'h1a7654c882c3e568;
    assign coff[7698] = 64'hba28423794bbe85a;
    assign coff[7699] = 64'h82c3e568e589ab38;
    assign coff[7700] = 64'h7d3c1a98e589ab38;
    assign coff[7701] = 64'h45d7bdc994bbe85a;
    assign coff[7702] = 64'he589ab3882c3e568;
    assign coff[7703] = 64'h94bbe85aba284237;
    assign coff[7704] = 64'h7dd4191de885cb9a;
    assign coff[7705] = 64'h485f8959966cc022;
    assign coff[7706] = 64'he885cb9a822be6e3;
    assign coff[7707] = 64'h966cc022b7a076a7;
    assign coff[7708] = 64'h69933fdeb7a076a7;
    assign coff[7709] = 64'h177a3466822be6e3;
    assign coff[7710] = 64'hb7a076a7966cc022;
    assign coff[7711] = 64'h822be6e3e885cb9a;
    assign coff[7712] = 64'h63e757eaaffacb76;
    assign coff[7713] = 64'h0e0f456f80c64612;
    assign coff[7714] = 64'haffacb769c18a816;
    assign coff[7715] = 64'h80c64612f1f0ba91;
    assign coff[7716] = 64'h7f39b9eef1f0ba91;
    assign coff[7717] = 64'h5005348a9c18a816;
    assign coff[7718] = 64'hf1f0ba9180c64612;
    assign coff[7719] = 64'h9c18a816affacb76;
    assign coff[7720] = 64'h7aebe28ddc4d65fb;
    assign coff[7721] = 64'h3dad300b8fd6e0c2;
    assign coff[7722] = 64'hdc4d65fb85141d73;
    assign coff[7723] = 64'h8fd6e0c2c252cff5;
    assign coff[7724] = 64'h70291f3ec252cff5;
    assign coff[7725] = 64'h23b29a0585141d73;
    assign coff[7726] = 64'hc252cff58fd6e0c2;
    assign coff[7727] = 64'h85141d73dc4d65fb;
    assign coff[7728] = 64'h719862b9c501ea0a;
    assign coff[7729] = 64'h269c268f85f6465c;
    assign coff[7730] = 64'hc501ea0a8e679d47;
    assign coff[7731] = 64'h85f6465cd963d971;
    assign coff[7732] = 64'h7a09b9a4d963d971;
    assign coff[7733] = 64'h3afe15f68e679d47;
    assign coff[7734] = 64'hd963d97185f6465c;
    assign coff[7735] = 64'h8e679d47c501ea0a;
    assign coff[7736] = 64'h7f861753f4f812e7;
    assign coff[7737] = 64'h525f74809e06e907;
    assign coff[7738] = 64'hf4f812e78079e8ad;
    assign coff[7739] = 64'h9e06e907ada08b80;
    assign coff[7740] = 64'h61f916f9ada08b80;
    assign coff[7741] = 64'h0b07ed198079e8ad;
    assign coff[7742] = 64'hada08b809e06e907;
    assign coff[7743] = 64'h8079e8adf4f812e7;
    assign coff[7744] = 64'h5fdb601bab2c8c27;
    assign coff[7745] = 64'h07ccd0a5803ce5c3;
    assign coff[7746] = 64'hab2c8c27a0249fe5;
    assign coff[7747] = 64'h803ce5c3f8332f5b;
    assign coff[7748] = 64'h7fc31a3df8332f5b;
    assign coff[7749] = 64'h54d373d9a0249fe5;
    assign coff[7750] = 64'hf8332f5b803ce5c3;
    assign coff[7751] = 64'ha0249fe5ab2c8c27;
    assign coff[7752] = 64'h79059212d65059ac;
    assign coff[7753] = 64'h381948648cf2b9b8;
    assign coff[7754] = 64'hd65059ac86fa6dee;
    assign coff[7755] = 64'h8cf2b9b8c7e6b79c;
    assign coff[7756] = 64'h730d4648c7e6b79c;
    assign coff[7757] = 64'h29afa65486fa6dee;
    assign coff[7758] = 64'hc7e6b79c8cf2b9b8;
    assign coff[7759] = 64'h86fa6deed65059ac;
    assign coff[7760] = 64'h6e905534bf8132ce;
    assign coff[7761] = 64'h209349338436ea23;
    assign coff[7762] = 64'hbf8132ce916faacc;
    assign coff[7763] = 64'h8436ea23df6cb6cd;
    assign coff[7764] = 64'h7bc915dddf6cb6cd;
    assign coff[7765] = 64'h407ecd32916faacc;
    assign coff[7766] = 64'hdf6cb6cd8436ea23;
    assign coff[7767] = 64'h916faaccbf8132ce;
    assign coff[7768] = 64'h7ed43438eeb99b8d;
    assign coff[7769] = 64'h4d7762319a1a68be;
    assign coff[7770] = 64'heeb99b8d812bcbc8;
    assign coff[7771] = 64'h9a1a68beb2889dcf;
    assign coff[7772] = 64'h65e59742b2889dcf;
    assign coff[7773] = 64'h11466473812bcbc8;
    assign coff[7774] = 64'hb2889dcf9a1a68be;
    assign coff[7775] = 64'h812bcbc8eeb99b8d;
    assign coff[7776] = 64'h67b5b2bbb4fa6489;
    assign coff[7777] = 64'h14490e74819e1cfd;
    assign coff[7778] = 64'hb4fa6489984a4d45;
    assign coff[7779] = 64'h819e1cfdebb6f18c;
    assign coff[7780] = 64'h7e61e303ebb6f18c;
    assign coff[7781] = 64'h4b059b77984a4d45;
    assign coff[7782] = 64'hebb6f18c819e1cfd;
    assign coff[7783] = 64'h984a4d45b4fa6489;
    assign coff[7784] = 64'h7c8663f4e260764f;
    assign coff[7785] = 64'h431b0e15930033f1;
    assign coff[7786] = 64'he260764f83799c0c;
    assign coff[7787] = 64'h930033f1bce4f1eb;
    assign coff[7788] = 64'h6cffcc0fbce4f1eb;
    assign coff[7789] = 64'h1d9f89b183799c0c;
    assign coff[7790] = 64'hbce4f1eb930033f1;
    assign coff[7791] = 64'h83799c0ce260764f;
    assign coff[7792] = 64'h745a619bcaa70322;
    assign coff[7793] = 64'h2c8d341a8800e62f;
    assign coff[7794] = 64'hcaa703228ba59e65;
    assign coff[7795] = 64'h8800e62fd372cbe6;
    assign coff[7796] = 64'h77ff19d1d372cbe6;
    assign coff[7797] = 64'h3558fcde8ba59e65;
    assign coff[7798] = 64'hd372cbe68800e62f;
    assign coff[7799] = 64'h8ba59e65caa70322;
    assign coff[7800] = 64'h7fe954bafb3d57d9;
    assign coff[7801] = 64'h5714b99da22fd57b;
    assign coff[7802] = 64'hfb3d57d98016ab46;
    assign coff[7803] = 64'ha22fd57ba8eb4663;
    assign coff[7804] = 64'h5dd02a85a8eb4663;
    assign coff[7805] = 64'h04c2a8278016ab46;
    assign coff[7806] = 64'ha8eb4663a22fd57b;
    assign coff[7807] = 64'h8016ab46fb3d57d9;
    assign coff[7808] = 64'h5dbf0f8ca8d8dc81;
    assign coff[7809] = 64'h04a98a888015be75;
    assign coff[7810] = 64'ha8d8dc81a240f074;
    assign coff[7811] = 64'h8015be75fb567578;
    assign coff[7812] = 64'h7fea418bfb567578;
    assign coff[7813] = 64'h5727237fa240f074;
    assign coff[7814] = 64'hfb5675788015be75;
    assign coff[7815] = 64'ha240f074a8d8dc81;
    assign coff[7816] = 64'h77f65819d35b3d13;
    assign coff[7817] = 64'h3542234c8b9b2718;
    assign coff[7818] = 64'hd35b3d138809a7e7;
    assign coff[7819] = 64'h8b9b2718cabddcb4;
    assign coff[7820] = 64'h7464d8e8cabddcb4;
    assign coff[7821] = 64'h2ca4c2ed8809a7e7;
    assign coff[7822] = 64'hcabddcb48b9b2718;
    assign coff[7823] = 64'h8809a7e7d35b3d13;
    assign coff[7824] = 64'h6cf29cdcbccf8c50;
    assign coff[7825] = 64'h1d8715d08373cd6c;
    assign coff[7826] = 64'hbccf8c50930d6324;
    assign coff[7827] = 64'h8373cd6ce278ea30;
    assign coff[7828] = 64'h7c8c3294e278ea30;
    assign coff[7829] = 64'h433073b0930d6324;
    assign coff[7830] = 64'he278ea308373cd6c;
    assign coff[7831] = 64'h930d6324bccf8c50;
    assign coff[7832] = 64'h7e5de4eceb9e2144;
    assign coff[7833] = 64'h4af13d00983b9442;
    assign coff[7834] = 64'heb9e214481a21b14;
    assign coff[7835] = 64'h983b9442b50ec300;
    assign coff[7836] = 64'h67c46bbeb50ec300;
    assign coff[7837] = 64'h1461debc81a21b14;
    assign coff[7838] = 64'hb50ec300983b9442;
    assign coff[7839] = 64'h81a21b14eb9e2144;
    assign coff[7840] = 64'h65d65f69b2749d68;
    assign coff[7841] = 64'h112d7d00812869e4;
    assign coff[7842] = 64'hb2749d689a29a097;
    assign coff[7843] = 64'h812869e4eed28300;
    assign coff[7844] = 64'h7ed7961ceed28300;
    assign coff[7845] = 64'h4d8b62989a29a097;
    assign coff[7846] = 64'heed28300812869e4;
    assign coff[7847] = 64'h9a29a097b2749d68;
    assign coff[7848] = 64'h7bc2ae10df54694b;
    assign coff[7849] = 64'h406916699163030b;
    assign coff[7850] = 64'hdf54694b843d51f0;
    assign coff[7851] = 64'h9163030bbf96e997;
    assign coff[7852] = 64'h6e9cfcf5bf96e997;
    assign coff[7853] = 64'h20ab96b5843d51f0;
    assign coff[7854] = 64'hbf96e9979163030b;
    assign coff[7855] = 64'h843d51f0df54694b;
    assign coff[7856] = 64'h7302403cc7d0218e;
    assign coff[7857] = 64'h2997e24f86f240e3;
    assign coff[7858] = 64'hc7d0218e8cfdbfc4;
    assign coff[7859] = 64'h86f240e3d6681db1;
    assign coff[7860] = 64'h790dbf1dd6681db1;
    assign coff[7861] = 64'h382fde728cfdbfc4;
    assign coff[7862] = 64'hd6681db186f240e3;
    assign coff[7863] = 64'h8cfdbfc4c7d0218e;
    assign coff[7864] = 64'h7fc18fb4f81a197b;
    assign coff[7865] = 64'h54c09feba013f9ed;
    assign coff[7866] = 64'hf81a197b803e704c;
    assign coff[7867] = 64'ha013f9edab3f6015;
    assign coff[7868] = 64'h5fec0613ab3f6015;
    assign coff[7869] = 64'h07e5e685803e704c;
    assign coff[7870] = 64'hab3f6015a013f9ed;
    assign coff[7871] = 64'h803e704cf81a197b;
    assign coff[7872] = 64'h61e8e893ad8d506e;
    assign coff[7873] = 64'h0aeee2d78077c0a8;
    assign coff[7874] = 64'had8d506e9e17176d;
    assign coff[7875] = 64'h8077c0a8f5111d29;
    assign coff[7876] = 64'h7f883f58f5111d29;
    assign coff[7877] = 64'h5272af929e17176d;
    assign coff[7878] = 64'hf5111d298077c0a8;
    assign coff[7879] = 64'h9e17176dad8d506e;
    assign coff[7880] = 64'h7a02228ad94be3e3;
    assign coff[7881] = 64'h3ae7c6e78e5c0a2e;
    assign coff[7882] = 64'hd94be3e385fddd76;
    assign coff[7883] = 64'h8e5c0a2ec5183919;
    assign coff[7884] = 64'h71a3f5d2c5183919;
    assign coff[7885] = 64'h26b41c1d85fddd76;
    assign coff[7886] = 64'hc51839198e5c0a2e;
    assign coff[7887] = 64'h85fddd76d94be3e3;
    assign coff[7888] = 64'h701d00e1c23ccb57;
    assign coff[7889] = 64'h239a76a0850d1d75;
    assign coff[7890] = 64'hc23ccb578fe2ff1f;
    assign coff[7891] = 64'h850d1d75dc658960;
    assign coff[7892] = 64'h7af2e28bdc658960;
    assign coff[7893] = 64'h3dc334a98fe2ff1f;
    assign coff[7894] = 64'hdc658960850d1d75;
    assign coff[7895] = 64'h8fe2ff1fc23ccb57;
    assign coff[7896] = 64'h7f36f4c3f1d7bfca;
    assign coff[7897] = 64'h4ff1954b9c08f3c1;
    assign coff[7898] = 64'hf1d7bfca80c90b3d;
    assign coff[7899] = 64'h9c08f3c1b00e6ab5;
    assign coff[7900] = 64'h63f70c3fb00e6ab5;
    assign coff[7901] = 64'h0e28403680c90b3d;
    assign coff[7902] = 64'hb00e6ab59c08f3c1;
    assign coff[7903] = 64'h80c90b3df1d7bfca;
    assign coff[7904] = 64'h698507f6b78bbd42;
    assign coff[7905] = 64'h17617f1d82274d36;
    assign coff[7906] = 64'hb78bbd42967af80a;
    assign coff[7907] = 64'h82274d36e89e80e3;
    assign coff[7908] = 64'h7dd8b2cae89e80e3;
    assign coff[7909] = 64'h487442be967af80a;
    assign coff[7910] = 64'he89e80e382274d36;
    assign coff[7911] = 64'h967af80ab78bbd42;
    assign coff[7912] = 64'h7d36e60be57114be;
    assign coff[7913] = 64'h45c2acaa94ae33be;
    assign coff[7914] = 64'he57114be82c919f5;
    assign coff[7915] = 64'h94ae33beba3d5356;
    assign coff[7916] = 64'h6b51cc42ba3d5356;
    assign coff[7917] = 64'h1a8eeb4282c919f5;
    assign coff[7918] = 64'hba3d535694ae33be;
    assign coff[7919] = 64'h82c919f5e57114be;
    assign coff[7920] = 64'h75a091c6cd861eaf;
    assign coff[7921] = 64'h2f7ba72989220c84;
    assign coff[7922] = 64'hcd861eaf8a5f6e3a;
    assign coff[7923] = 64'h89220c84d08458d7;
    assign coff[7924] = 64'h76ddf37cd08458d7;
    assign coff[7925] = 64'h3279e1518a5f6e3a;
    assign coff[7926] = 64'hd08458d789220c84;
    assign coff[7927] = 64'h8a5f6e3acd861eaf;
    assign coff[7928] = 64'h7ffd6042fe615223;
    assign coff[7929] = 64'h595b65aaa45a2872;
    assign coff[7930] = 64'hfe61522380029fbe;
    assign coff[7931] = 64'ha45a2872a6a49a56;
    assign coff[7932] = 64'h5ba5d78ea6a49a56;
    assign coff[7933] = 64'h019eaddd80029fbe;
    assign coff[7934] = 64'ha6a49a56a45a2872;
    assign coff[7935] = 64'h80029fbefe615223;
    assign coff[7936] = 64'h5cab762fa7b40933;
    assign coff[7937] = 64'h03179ab580099029;
    assign coff[7938] = 64'ha7b40933a35489d1;
    assign coff[7939] = 64'h80099029fce8654b;
    assign coff[7940] = 64'h7ff66fd7fce8654b;
    assign coff[7941] = 64'h584bf6cda35489d1;
    assign coff[7942] = 64'hfce8654b80099029;
    assign coff[7943] = 64'ha35489d1a7b40933;
    assign coff[7944] = 64'h7767c880d1e33c69;
    assign coff[7945] = 64'h33d375468af615a3;
    assign coff[7946] = 64'hd1e33c6988983780;
    assign coff[7947] = 64'h8af615a3cc2c8aba;
    assign coff[7948] = 64'h7509ea5dcc2c8aba;
    assign coff[7949] = 64'h2e1cc39788983780;
    assign coff[7950] = 64'hcc2c8aba8af615a3;
    assign coff[7951] = 64'h88983780d1e33c69;
    assign coff[7952] = 64'h6c1d6fc6bb7a9521;
    assign coff[7953] = 64'h1bff3f7583197110;
    assign coff[7954] = 64'hbb7a952193e2903a;
    assign coff[7955] = 64'h83197110e400c08b;
    assign coff[7956] = 64'h7ce68ef0e400c08b;
    assign coff[7957] = 64'h44856adf93e2903a;
    assign coff[7958] = 64'he400c08b83197110;
    assign coff[7959] = 64'h93e2903abb7a9521;
    assign coff[7960] = 64'h7e1b6d53ea118a35;
    assign coff[7961] = 64'h49a9ceaf975225a1;
    assign coff[7962] = 64'hea118a3581e492ad;
    assign coff[7963] = 64'h975225a1b6563151;
    assign coff[7964] = 64'h68adda5fb6563151;
    assign coff[7965] = 64'h15ee75cb81e492ad;
    assign coff[7966] = 64'hb6563151975225a1;
    assign coff[7967] = 64'h81e492adea118a35;
    assign coff[7968] = 64'h64e0cd78b1362fa2;
    assign coff[7969] = 64'h0f9eae4c80f4e50e;
    assign coff[7970] = 64'hb1362fa29b1f3288;
    assign coff[7971] = 64'h80f4e50ef06151b4;
    assign coff[7972] = 64'h7f0b1af2f06151b4;
    assign coff[7973] = 64'h4ec9d05e9b1f3288;
    assign coff[7974] = 64'hf06151b480f4e50e;
    assign coff[7975] = 64'h9b1f3288b1362fa2;
    assign coff[7976] = 64'h7b59a902ddd03eef;
    assign coff[7977] = 64'h3f0c5a5a909acc32;
    assign coff[7978] = 64'hddd03eef84a656fe;
    assign coff[7979] = 64'h909acc32c0f3a5a6;
    assign coff[7980] = 64'h6f6533cec0f3a5a6;
    assign coff[7981] = 64'h222fc11184a656fe;
    assign coff[7982] = 64'hc0f3a5a6909acc32;
    assign coff[7983] = 64'h84a656feddd03eef;
    assign coff[7984] = 64'h724f8593c667e996;
    assign coff[7985] = 64'h281aca578671ebc8;
    assign coff[7986] = 64'hc667e9968db07a6d;
    assign coff[7987] = 64'h8671ebc8d7e535a9;
    assign coff[7988] = 64'h798e1438d7e535a9;
    assign coff[7989] = 64'h3998166a8db07a6d;
    assign coff[7990] = 64'hd7e535a98671ebc8;
    assign coff[7991] = 64'h8db07a6dc667e996;
    assign coff[7992] = 64'h7fa6496ef688e77c;
    assign coff[7993] = 64'h5391a6999f0b9307;
    assign coff[7994] = 64'hf688e77c8059b692;
    assign coff[7995] = 64'h9f0b9307ac6e5967;
    assign coff[7996] = 64'h60f46cf9ac6e5967;
    assign coff[7997] = 64'h097718848059b692;
    assign coff[7998] = 64'hac6e59679f0b9307;
    assign coff[7999] = 64'h8059b692f688e77c;
    assign coff[8000] = 64'h60e40278ac5b5189;
    assign coff[8001] = 64'h095e07f88057dd41;
    assign coff[8002] = 64'hac5b51899f1bfd88;
    assign coff[8003] = 64'h8057dd41f6a1f808;
    assign coff[8004] = 64'h7fa822bff6a1f808;
    assign coff[8005] = 64'h53a4ae779f1bfd88;
    assign coff[8006] = 64'hf6a1f8088057dd41;
    assign coff[8007] = 64'h9f1bfd88ac5b5189;
    assign coff[8008] = 64'h798631ffd7cd586a;
    assign coff[8009] = 64'h3981a36d8da52da3;
    assign coff[8010] = 64'hd7cd586a8679ce01;
    assign coff[8011] = 64'h8da52da3c67e5c93;
    assign coff[8012] = 64'h725ad25dc67e5c93;
    assign coff[8013] = 64'h2832a7968679ce01;
    assign coff[8014] = 64'hc67e5c938da52da3;
    assign coff[8015] = 64'h8679ce01d7cd586a;
    assign coff[8016] = 64'h6f58d082c0ddc786;
    assign coff[8017] = 64'h22178826849fa2f7;
    assign coff[8018] = 64'hc0ddc78690a72f7e;
    assign coff[8019] = 64'h849fa2f7dde877da;
    assign coff[8020] = 64'h7b605d09dde877da;
    assign coff[8021] = 64'h3f22387a90a72f7e;
    assign coff[8022] = 64'hdde877da849fa2f7;
    assign coff[8023] = 64'h90a72f7ec0ddc786;
    assign coff[8024] = 64'h7f08075cf048601c;
    assign coff[8025] = 64'h4eb600299b0fbc24;
    assign coff[8026] = 64'hf048601c80f7f8a4;
    assign coff[8027] = 64'h9b0fbc24b149ffd7;
    assign coff[8028] = 64'h64f043dcb149ffd7;
    assign coff[8029] = 64'h0fb79fe480f7f8a4;
    assign coff[8030] = 64'hb149ffd79b0fbc24;
    assign coff[8031] = 64'h80f7f8a4f048601c;
    assign coff[8032] = 64'h689f61a1b641a4fe;
    assign coff[8033] = 64'h15d5b28881e046b6;
    assign coff[8034] = 64'hb641a4fe97609e5f;
    assign coff[8035] = 64'h81e046b6ea2a4d78;
    assign coff[8036] = 64'h7e1fb94aea2a4d78;
    assign coff[8037] = 64'h49be5b0297609e5f;
    assign coff[8038] = 64'hea2a4d7881e046b6;
    assign coff[8039] = 64'h97609e5fb641a4fe;
    assign coff[8040] = 64'h7ce10d3fe3e83ae5;
    assign coff[8041] = 64'h44702f1993d51e10;
    assign coff[8042] = 64'he3e83ae5831ef2c1;
    assign coff[8043] = 64'h93d51e10bb8fd0e7;
    assign coff[8044] = 64'h6c2ae1f0bb8fd0e7;
    assign coff[8045] = 64'h1c17c51b831ef2c1;
    assign coff[8046] = 64'hbb8fd0e793d51e10;
    assign coff[8047] = 64'h831ef2c1e3e83ae5;
    assign coff[8048] = 64'h74ffbb0dcc1590b8;
    assign coff[8049] = 64'h2e0550bb888f2bf1;
    assign coff[8050] = 64'hcc1590b88b0044f3;
    assign coff[8051] = 64'h888f2bf1d1faaf45;
    assign coff[8052] = 64'h7770d40fd1faaf45;
    assign coff[8053] = 64'h33ea6f488b0044f3;
    assign coff[8054] = 64'hd1faaf45888f2bf1;
    assign coff[8055] = 64'h8b0044f3cc1590b8;
    assign coff[8056] = 64'h7ff5d1f1fccf453f;
    assign coff[8057] = 64'h5839c302a3433554;
    assign coff[8058] = 64'hfccf453f800a2e0f;
    assign coff[8059] = 64'ha3433554a7c63cfe;
    assign coff[8060] = 64'h5cbccaaca7c63cfe;
    assign coff[8061] = 64'h0330bac1800a2e0f;
    assign coff[8062] = 64'ha7c63cfea3433554;
    assign coff[8063] = 64'h800a2e0ffccf453f;
    assign coff[8064] = 64'h5ecf0bafaa010bf6;
    assign coff[8065] = 64'h063b4c578026db36;
    assign coff[8066] = 64'haa010bf6a130f451;
    assign coff[8067] = 64'h8026db36f9c4b3a9;
    assign coff[8068] = 64'h7fd924caf9c4b3a9;
    assign coff[8069] = 64'h55fef40aa130f451;
    assign coff[8070] = 64'hf9c4b3a98026db36;
    assign coff[8071] = 64'ha130f451aa010bf6;
    assign coff[8072] = 64'h788047bad4d4f65a;
    assign coff[8073] = 64'h36aec3b08c44b54d;
    assign coff[8074] = 64'hd4d4f65a877fb846;
    assign coff[8075] = 64'h8c44b54dc9513c50;
    assign coff[8076] = 64'h73bb4ab3c9513c50;
    assign coff[8077] = 64'h2b2b09a6877fb846;
    assign coff[8078] = 64'hc9513c508c44b54d;
    assign coff[8079] = 64'h877fb846d4d4f65a;
    assign coff[8080] = 64'h6dc396b0be271a9f;
    assign coff[8081] = 64'h1f0dc8c083d2f701;
    assign coff[8082] = 64'hbe271a9f923c6950;
    assign coff[8083] = 64'h83d2f701e0f23740;
    assign coff[8084] = 64'h7c2d08ffe0f23740;
    assign coff[8085] = 64'h41d8e561923c6950;
    assign coff[8086] = 64'he0f2374083d2f701;
    assign coff[8087] = 64'h923c6950be271a9f;
    assign coff[8088] = 64'h7e9b7d58ed2b817d;
    assign coff[8089] = 64'h4c35c7ac99290303;
    assign coff[8090] = 64'hed2b817d816482a8;
    assign coff[8091] = 64'h99290303b3ca3854;
    assign coff[8092] = 64'h66d6fcfdb3ca3854;
    assign coff[8093] = 64'h12d47e83816482a8;
    assign coff[8094] = 64'hb3ca385499290303;
    assign coff[8095] = 64'h816482a8ed2b817d;
    assign coff[8096] = 64'h66c80445b3b60881;
    assign coff[8097] = 64'h12bba22b8160d298;
    assign coff[8098] = 64'hb3b608819937fbbb;
    assign coff[8099] = 64'h8160d298ed445dd5;
    assign coff[8100] = 64'h7e9f2d68ed445dd5;
    assign coff[8101] = 64'h4c49f77f9937fbbb;
    assign coff[8102] = 64'hed445dd58160d298;
    assign coff[8103] = 64'h9937fbbbb3b60881;
    assign coff[8104] = 64'h7c26edabe0d9d616;
    assign coff[8105] = 64'h41c356c5922f7d96;
    assign coff[8106] = 64'he0d9d61683d91255;
    assign coff[8107] = 64'h922f7d96be3ca93b;
    assign coff[8108] = 64'h6dd0826abe3ca93b;
    assign coff[8109] = 64'h1f2629ea83d91255;
    assign coff[8110] = 64'hbe3ca93b922f7d96;
    assign coff[8111] = 64'h83d91255e0d9d616;
    assign coff[8112] = 64'h73b08bd1c93a8410;
    assign coff[8113] = 64'h2b135fc6877740bb;
    assign coff[8114] = 64'hc93a84108c4f742f;
    assign coff[8115] = 64'h877740bbd4eca03a;
    assign coff[8116] = 64'h7888bf45d4eca03a;
    assign coff[8117] = 64'h36c57bf08c4f742f;
    assign coff[8118] = 64'hd4eca03a877740bb;
    assign coff[8119] = 64'h8c4f742fc93a8410;
    assign coff[8120] = 64'h7fd7e917f9ab996e;
    assign coff[8121] = 64'h55ec54c6a1201385;
    assign coff[8122] = 64'hf9ab996e802816e9;
    assign coff[8123] = 64'ha1201385aa13ab3a;
    assign coff[8124] = 64'h5edfec7baa13ab3a;
    assign coff[8125] = 64'h06546692802816e9;
    assign coff[8126] = 64'haa13ab3aa1201385;
    assign coff[8127] = 64'h802816e9f9ab996e;
    assign coff[8128] = 64'h62ea085caec27d0c;
    assign coff[8129] = 64'h0c7f51cf809c8ebc;
    assign coff[8130] = 64'haec27d0c9d15f7a4;
    assign coff[8131] = 64'h809c8ebcf380ae31;
    assign coff[8132] = 64'h7f637144f380ae31;
    assign coff[8133] = 64'h513d82f49d15f7a4;
    assign coff[8134] = 64'hf380ae31809c8ebc;
    assign coff[8135] = 64'h9d15f7a4aec27d0c;
    assign coff[8136] = 64'h7a795eecdacbed58;
    assign coff[8137] = 64'h3c4ba5048f17484b;
    assign coff[8138] = 64'hdacbed588586a114;
    assign coff[8139] = 64'h8f17484bc3b45afc;
    assign coff[8140] = 64'h70e8b7b5c3b45afc;
    assign coff[8141] = 64'h253412a88586a114;
    assign coff[8142] = 64'hc3b45afc8f17484b;
    assign coff[8143] = 64'h8586a114dacbed58;
    assign coff[8144] = 64'h70dcdec0c39e30b8;
    assign coff[8145] = 64'h251c05b8857f5564;
    assign coff[8146] = 64'hc39e30b88f232140;
    assign coff[8147] = 64'h857f5564dae3fa48;
    assign coff[8148] = 64'h7a80aa9cdae3fa48;
    assign coff[8149] = 64'h3c61cf488f232140;
    assign coff[8150] = 64'hdae3fa48857f5564;
    assign coff[8151] = 64'h8f232140c39e30b8;
    assign coff[8152] = 64'h7f60faa0f367ab31;
    assign coff[8153] = 64'h512a156b9d0605f7;
    assign coff[8154] = 64'hf367ab31809f0560;
    assign coff[8155] = 64'h9d0605f7aed5ea95;
    assign coff[8156] = 64'h62f9fa09aed5ea95;
    assign coff[8157] = 64'h0c9854cf809f0560;
    assign coff[8158] = 64'haed5ea959d0605f7;
    assign coff[8159] = 64'h809f0560f367ab31;
    assign coff[8160] = 64'h6a669cddb8d8a09d;
    assign coff[8161] = 64'h18ec64f082732dc0;
    assign coff[8162] = 64'hb8d8a09d95996323;
    assign coff[8163] = 64'h82732dc0e7139b10;
    assign coff[8164] = 64'h7d8cd240e7139b10;
    assign coff[8165] = 64'h47275f6395996323;
    assign coff[8166] = 64'he7139b1082732dc0;
    assign coff[8167] = 64'h95996323b8d8a09d;
    assign coff[8168] = 64'h7d87eb0ae6faf4b5;
    assign coff[8169] = 64'h471279ba958b6c9b;
    assign coff[8170] = 64'he6faf4b5827814f6;
    assign coff[8171] = 64'h958b6c9bb8ed8646;
    assign coff[8172] = 64'h6a749365b8ed8646;
    assign coff[8173] = 64'h19050b4b827814f6;
    assign coff[8174] = 64'hb8ed8646958b6c9b;
    assign coff[8175] = 64'h827814f6e6faf4b5;
    assign coff[8176] = 64'h763cdf94cef89ed2;
    assign coff[8177] = 64'h30f028f489b9823e;
    assign coff[8178] = 64'hcef89ed289c3206c;
    assign coff[8179] = 64'h89b9823ecf0fd70c;
    assign coff[8180] = 64'h76467dc2cf0fd70c;
    assign coff[8181] = 64'h3107612e89c3206c;
    assign coff[8182] = 64'hcf0fd70c89b9823e;
    assign coff[8183] = 64'h89c3206ccef89ed2;
    assign coff[8184] = 64'h7fffff62fff36f02;
    assign coff[8185] = 64'h5a799669a574a414;
    assign coff[8186] = 64'hfff36f028000009e;
    assign coff[8187] = 64'ha574a414a5866997;
    assign coff[8188] = 64'h5a8b5beca5866997;
    assign coff[8189] = 64'h000c90fe8000009e;
    assign coff[8190] = 64'ha5866997a574a414;
    assign coff[8191] = 64'h8000009efff36f02;

    always_ff @(posedge clk, negedge rst_n) begin
        if(~rst_n) begin
            data_o <= 'b0;
        end else begin
            data_o <= coff[addr_i];
        end
    end

endmodule